module main (input  I0, input  I1, output  O);
wire  inst0_0;
xor inst0 (inst0_0, I0, I1);
assign O = inst0_0;
endmodule

