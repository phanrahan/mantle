module Or4x8 (
    input [7:0] I0,
    input [7:0] I1,
    input [7:0] I2,
    input [7:0] I3,
    output [7:0] O
);
assign O = {| ({I3[7],I2[7],I1[7],I0[7]}),| ({I3[6],I2[6],I1[6],I0[6]}),| ({I3[5],I2[5],I1[5],I0[5]}),| ({I3[4],I2[4],I1[4],I0[4]}),| ({I3[3],I2[3],I1[3],I0[3]}),| ({I3[2],I2[2],I1[2],I0[2]}),| ({I3[1],I2[1],I1[1],I0[1]}),| ({I3[0],I2[0],I1[0],I0[0]})};
endmodule

