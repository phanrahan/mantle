module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk, input [width-1:0] in, output [width-1:0] out);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse (input I, output O, input CLK);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1'b1), .init(1'h1), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input I, output O, input CLK);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1'b1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Ring8_0001 (output [7:0] O, input CLK);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.I(DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O), .CLK(CLK));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O), .CLK(CLK));
DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.I(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O), .O(DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O), .CLK(CLK));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O,DFF_init1_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

