module Decode_0_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0001)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_1_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0002)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_2_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0004)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_3_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0008)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_4_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0010)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_5_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0020)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_6_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0040)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_7_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0080)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_8_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0100)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_9_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0200)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_10_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0400)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_11_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0800)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_12_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h1000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_13_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h2000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_14_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h4000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_15_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h8000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_16_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_17_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_18_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_19_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_20_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_21_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_22_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_23_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_24_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_25_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_26_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_27_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_28_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_29_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_30_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_31_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_32_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_33_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_34_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_35_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_36_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_37_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_38_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_39_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_40_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_41_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_42_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_43_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_44_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_45_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_46_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_47_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_48_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_49_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_50_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_51_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_52_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_53_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_54_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_55_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_56_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_57_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_58_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_59_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_60_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_61_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_62_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_63_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_64_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_65_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_66_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_67_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_68_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_69_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_70_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_71_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_72_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_73_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_74_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_75_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_76_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_77_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_78_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_79_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_80_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_81_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_82_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_83_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_84_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_85_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_86_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_87_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_88_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_89_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_90_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_91_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_92_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_93_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_94_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_95_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_96_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_97_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_98_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_99_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_100_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_101_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_102_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_103_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_104_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_105_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_106_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_107_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_108_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_109_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_110_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_111_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_112_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_113_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_114_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_115_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_116_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_117_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_118_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_119_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_120_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_121_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_122_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_123_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_124_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_125_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_126_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_127_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_128_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_129_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_130_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_131_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_132_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_133_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_134_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_135_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_136_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_137_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_138_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_139_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_140_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_141_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_142_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_143_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_144_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_145_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_146_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_147_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_148_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_149_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_150_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_151_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_152_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_153_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_154_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_155_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_156_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_157_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_158_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_159_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_160_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_161_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_162_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_163_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_164_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_165_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_166_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_167_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_168_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_169_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_170_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_171_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_172_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_173_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_174_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_175_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_176_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_177_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_178_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_179_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_180_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_181_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_182_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_183_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_184_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_185_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_186_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_187_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_188_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_189_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_190_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_191_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_192_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_193_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_194_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_195_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_196_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_197_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_198_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_199_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_200_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_201_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_202_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_203_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_204_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_205_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_206_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_207_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_208_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_209_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_210_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_211_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_212_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_213_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_214_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_215_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_216_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_217_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_218_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_219_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_220_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_221_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_222_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_223_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_224_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_225_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_226_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_227_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_228_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_229_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_230_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_231_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_232_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_233_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_234_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_235_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_236_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_237_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_238_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_239_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_240_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0001)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_241_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0002)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_242_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0004)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_243_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0008)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_244_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0010)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_245_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0020)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_246_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0040)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_247_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0080)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_248_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0100)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_249_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0200)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_250_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0400)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_251_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0800)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_252_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h1000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_253_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h2000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_254_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h4000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decode_255_8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0000)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h8000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire  Decode_0_8_inst0_O;
wire  Decode_1_8_inst0_O;
wire  Decode_2_8_inst0_O;
wire  Decode_3_8_inst0_O;
wire  Decode_4_8_inst0_O;
wire  Decode_5_8_inst0_O;
wire  Decode_6_8_inst0_O;
wire  Decode_7_8_inst0_O;
wire  Decode_8_8_inst0_O;
wire  Decode_9_8_inst0_O;
wire  Decode_10_8_inst0_O;
wire  Decode_11_8_inst0_O;
wire  Decode_12_8_inst0_O;
wire  Decode_13_8_inst0_O;
wire  Decode_14_8_inst0_O;
wire  Decode_15_8_inst0_O;
wire  Decode_16_8_inst0_O;
wire  Decode_17_8_inst0_O;
wire  Decode_18_8_inst0_O;
wire  Decode_19_8_inst0_O;
wire  Decode_20_8_inst0_O;
wire  Decode_21_8_inst0_O;
wire  Decode_22_8_inst0_O;
wire  Decode_23_8_inst0_O;
wire  Decode_24_8_inst0_O;
wire  Decode_25_8_inst0_O;
wire  Decode_26_8_inst0_O;
wire  Decode_27_8_inst0_O;
wire  Decode_28_8_inst0_O;
wire  Decode_29_8_inst0_O;
wire  Decode_30_8_inst0_O;
wire  Decode_31_8_inst0_O;
wire  Decode_32_8_inst0_O;
wire  Decode_33_8_inst0_O;
wire  Decode_34_8_inst0_O;
wire  Decode_35_8_inst0_O;
wire  Decode_36_8_inst0_O;
wire  Decode_37_8_inst0_O;
wire  Decode_38_8_inst0_O;
wire  Decode_39_8_inst0_O;
wire  Decode_40_8_inst0_O;
wire  Decode_41_8_inst0_O;
wire  Decode_42_8_inst0_O;
wire  Decode_43_8_inst0_O;
wire  Decode_44_8_inst0_O;
wire  Decode_45_8_inst0_O;
wire  Decode_46_8_inst0_O;
wire  Decode_47_8_inst0_O;
wire  Decode_48_8_inst0_O;
wire  Decode_49_8_inst0_O;
wire  Decode_50_8_inst0_O;
wire  Decode_51_8_inst0_O;
wire  Decode_52_8_inst0_O;
wire  Decode_53_8_inst0_O;
wire  Decode_54_8_inst0_O;
wire  Decode_55_8_inst0_O;
wire  Decode_56_8_inst0_O;
wire  Decode_57_8_inst0_O;
wire  Decode_58_8_inst0_O;
wire  Decode_59_8_inst0_O;
wire  Decode_60_8_inst0_O;
wire  Decode_61_8_inst0_O;
wire  Decode_62_8_inst0_O;
wire  Decode_63_8_inst0_O;
wire  Decode_64_8_inst0_O;
wire  Decode_65_8_inst0_O;
wire  Decode_66_8_inst0_O;
wire  Decode_67_8_inst0_O;
wire  Decode_68_8_inst0_O;
wire  Decode_69_8_inst0_O;
wire  Decode_70_8_inst0_O;
wire  Decode_71_8_inst0_O;
wire  Decode_72_8_inst0_O;
wire  Decode_73_8_inst0_O;
wire  Decode_74_8_inst0_O;
wire  Decode_75_8_inst0_O;
wire  Decode_76_8_inst0_O;
wire  Decode_77_8_inst0_O;
wire  Decode_78_8_inst0_O;
wire  Decode_79_8_inst0_O;
wire  Decode_80_8_inst0_O;
wire  Decode_81_8_inst0_O;
wire  Decode_82_8_inst0_O;
wire  Decode_83_8_inst0_O;
wire  Decode_84_8_inst0_O;
wire  Decode_85_8_inst0_O;
wire  Decode_86_8_inst0_O;
wire  Decode_87_8_inst0_O;
wire  Decode_88_8_inst0_O;
wire  Decode_89_8_inst0_O;
wire  Decode_90_8_inst0_O;
wire  Decode_91_8_inst0_O;
wire  Decode_92_8_inst0_O;
wire  Decode_93_8_inst0_O;
wire  Decode_94_8_inst0_O;
wire  Decode_95_8_inst0_O;
wire  Decode_96_8_inst0_O;
wire  Decode_97_8_inst0_O;
wire  Decode_98_8_inst0_O;
wire  Decode_99_8_inst0_O;
wire  Decode_100_8_inst0_O;
wire  Decode_101_8_inst0_O;
wire  Decode_102_8_inst0_O;
wire  Decode_103_8_inst0_O;
wire  Decode_104_8_inst0_O;
wire  Decode_105_8_inst0_O;
wire  Decode_106_8_inst0_O;
wire  Decode_107_8_inst0_O;
wire  Decode_108_8_inst0_O;
wire  Decode_109_8_inst0_O;
wire  Decode_110_8_inst0_O;
wire  Decode_111_8_inst0_O;
wire  Decode_112_8_inst0_O;
wire  Decode_113_8_inst0_O;
wire  Decode_114_8_inst0_O;
wire  Decode_115_8_inst0_O;
wire  Decode_116_8_inst0_O;
wire  Decode_117_8_inst0_O;
wire  Decode_118_8_inst0_O;
wire  Decode_119_8_inst0_O;
wire  Decode_120_8_inst0_O;
wire  Decode_121_8_inst0_O;
wire  Decode_122_8_inst0_O;
wire  Decode_123_8_inst0_O;
wire  Decode_124_8_inst0_O;
wire  Decode_125_8_inst0_O;
wire  Decode_126_8_inst0_O;
wire  Decode_127_8_inst0_O;
wire  Decode_128_8_inst0_O;
wire  Decode_129_8_inst0_O;
wire  Decode_130_8_inst0_O;
wire  Decode_131_8_inst0_O;
wire  Decode_132_8_inst0_O;
wire  Decode_133_8_inst0_O;
wire  Decode_134_8_inst0_O;
wire  Decode_135_8_inst0_O;
wire  Decode_136_8_inst0_O;
wire  Decode_137_8_inst0_O;
wire  Decode_138_8_inst0_O;
wire  Decode_139_8_inst0_O;
wire  Decode_140_8_inst0_O;
wire  Decode_141_8_inst0_O;
wire  Decode_142_8_inst0_O;
wire  Decode_143_8_inst0_O;
wire  Decode_144_8_inst0_O;
wire  Decode_145_8_inst0_O;
wire  Decode_146_8_inst0_O;
wire  Decode_147_8_inst0_O;
wire  Decode_148_8_inst0_O;
wire  Decode_149_8_inst0_O;
wire  Decode_150_8_inst0_O;
wire  Decode_151_8_inst0_O;
wire  Decode_152_8_inst0_O;
wire  Decode_153_8_inst0_O;
wire  Decode_154_8_inst0_O;
wire  Decode_155_8_inst0_O;
wire  Decode_156_8_inst0_O;
wire  Decode_157_8_inst0_O;
wire  Decode_158_8_inst0_O;
wire  Decode_159_8_inst0_O;
wire  Decode_160_8_inst0_O;
wire  Decode_161_8_inst0_O;
wire  Decode_162_8_inst0_O;
wire  Decode_163_8_inst0_O;
wire  Decode_164_8_inst0_O;
wire  Decode_165_8_inst0_O;
wire  Decode_166_8_inst0_O;
wire  Decode_167_8_inst0_O;
wire  Decode_168_8_inst0_O;
wire  Decode_169_8_inst0_O;
wire  Decode_170_8_inst0_O;
wire  Decode_171_8_inst0_O;
wire  Decode_172_8_inst0_O;
wire  Decode_173_8_inst0_O;
wire  Decode_174_8_inst0_O;
wire  Decode_175_8_inst0_O;
wire  Decode_176_8_inst0_O;
wire  Decode_177_8_inst0_O;
wire  Decode_178_8_inst0_O;
wire  Decode_179_8_inst0_O;
wire  Decode_180_8_inst0_O;
wire  Decode_181_8_inst0_O;
wire  Decode_182_8_inst0_O;
wire  Decode_183_8_inst0_O;
wire  Decode_184_8_inst0_O;
wire  Decode_185_8_inst0_O;
wire  Decode_186_8_inst0_O;
wire  Decode_187_8_inst0_O;
wire  Decode_188_8_inst0_O;
wire  Decode_189_8_inst0_O;
wire  Decode_190_8_inst0_O;
wire  Decode_191_8_inst0_O;
wire  Decode_192_8_inst0_O;
wire  Decode_193_8_inst0_O;
wire  Decode_194_8_inst0_O;
wire  Decode_195_8_inst0_O;
wire  Decode_196_8_inst0_O;
wire  Decode_197_8_inst0_O;
wire  Decode_198_8_inst0_O;
wire  Decode_199_8_inst0_O;
wire  Decode_200_8_inst0_O;
wire  Decode_201_8_inst0_O;
wire  Decode_202_8_inst0_O;
wire  Decode_203_8_inst0_O;
wire  Decode_204_8_inst0_O;
wire  Decode_205_8_inst0_O;
wire  Decode_206_8_inst0_O;
wire  Decode_207_8_inst0_O;
wire  Decode_208_8_inst0_O;
wire  Decode_209_8_inst0_O;
wire  Decode_210_8_inst0_O;
wire  Decode_211_8_inst0_O;
wire  Decode_212_8_inst0_O;
wire  Decode_213_8_inst0_O;
wire  Decode_214_8_inst0_O;
wire  Decode_215_8_inst0_O;
wire  Decode_216_8_inst0_O;
wire  Decode_217_8_inst0_O;
wire  Decode_218_8_inst0_O;
wire  Decode_219_8_inst0_O;
wire  Decode_220_8_inst0_O;
wire  Decode_221_8_inst0_O;
wire  Decode_222_8_inst0_O;
wire  Decode_223_8_inst0_O;
wire  Decode_224_8_inst0_O;
wire  Decode_225_8_inst0_O;
wire  Decode_226_8_inst0_O;
wire  Decode_227_8_inst0_O;
wire  Decode_228_8_inst0_O;
wire  Decode_229_8_inst0_O;
wire  Decode_230_8_inst0_O;
wire  Decode_231_8_inst0_O;
wire  Decode_232_8_inst0_O;
wire  Decode_233_8_inst0_O;
wire  Decode_234_8_inst0_O;
wire  Decode_235_8_inst0_O;
wire  Decode_236_8_inst0_O;
wire  Decode_237_8_inst0_O;
wire  Decode_238_8_inst0_O;
wire  Decode_239_8_inst0_O;
wire  Decode_240_8_inst0_O;
wire  Decode_241_8_inst0_O;
wire  Decode_242_8_inst0_O;
wire  Decode_243_8_inst0_O;
wire  Decode_244_8_inst0_O;
wire  Decode_245_8_inst0_O;
wire  Decode_246_8_inst0_O;
wire  Decode_247_8_inst0_O;
wire  Decode_248_8_inst0_O;
wire  Decode_249_8_inst0_O;
wire  Decode_250_8_inst0_O;
wire  Decode_251_8_inst0_O;
wire  Decode_252_8_inst0_O;
wire  Decode_253_8_inst0_O;
wire  Decode_254_8_inst0_O;
wire  Decode_255_8_inst0_O;
Decode_0_8 Decode_0_8_inst0 (.I(I), .O(Decode_0_8_inst0_O));
Decode_1_8 Decode_1_8_inst0 (.I(I), .O(Decode_1_8_inst0_O));
Decode_2_8 Decode_2_8_inst0 (.I(I), .O(Decode_2_8_inst0_O));
Decode_3_8 Decode_3_8_inst0 (.I(I), .O(Decode_3_8_inst0_O));
Decode_4_8 Decode_4_8_inst0 (.I(I), .O(Decode_4_8_inst0_O));
Decode_5_8 Decode_5_8_inst0 (.I(I), .O(Decode_5_8_inst0_O));
Decode_6_8 Decode_6_8_inst0 (.I(I), .O(Decode_6_8_inst0_O));
Decode_7_8 Decode_7_8_inst0 (.I(I), .O(Decode_7_8_inst0_O));
Decode_8_8 Decode_8_8_inst0 (.I(I), .O(Decode_8_8_inst0_O));
Decode_9_8 Decode_9_8_inst0 (.I(I), .O(Decode_9_8_inst0_O));
Decode_10_8 Decode_10_8_inst0 (.I(I), .O(Decode_10_8_inst0_O));
Decode_11_8 Decode_11_8_inst0 (.I(I), .O(Decode_11_8_inst0_O));
Decode_12_8 Decode_12_8_inst0 (.I(I), .O(Decode_12_8_inst0_O));
Decode_13_8 Decode_13_8_inst0 (.I(I), .O(Decode_13_8_inst0_O));
Decode_14_8 Decode_14_8_inst0 (.I(I), .O(Decode_14_8_inst0_O));
Decode_15_8 Decode_15_8_inst0 (.I(I), .O(Decode_15_8_inst0_O));
Decode_16_8 Decode_16_8_inst0 (.I(I), .O(Decode_16_8_inst0_O));
Decode_17_8 Decode_17_8_inst0 (.I(I), .O(Decode_17_8_inst0_O));
Decode_18_8 Decode_18_8_inst0 (.I(I), .O(Decode_18_8_inst0_O));
Decode_19_8 Decode_19_8_inst0 (.I(I), .O(Decode_19_8_inst0_O));
Decode_20_8 Decode_20_8_inst0 (.I(I), .O(Decode_20_8_inst0_O));
Decode_21_8 Decode_21_8_inst0 (.I(I), .O(Decode_21_8_inst0_O));
Decode_22_8 Decode_22_8_inst0 (.I(I), .O(Decode_22_8_inst0_O));
Decode_23_8 Decode_23_8_inst0 (.I(I), .O(Decode_23_8_inst0_O));
Decode_24_8 Decode_24_8_inst0 (.I(I), .O(Decode_24_8_inst0_O));
Decode_25_8 Decode_25_8_inst0 (.I(I), .O(Decode_25_8_inst0_O));
Decode_26_8 Decode_26_8_inst0 (.I(I), .O(Decode_26_8_inst0_O));
Decode_27_8 Decode_27_8_inst0 (.I(I), .O(Decode_27_8_inst0_O));
Decode_28_8 Decode_28_8_inst0 (.I(I), .O(Decode_28_8_inst0_O));
Decode_29_8 Decode_29_8_inst0 (.I(I), .O(Decode_29_8_inst0_O));
Decode_30_8 Decode_30_8_inst0 (.I(I), .O(Decode_30_8_inst0_O));
Decode_31_8 Decode_31_8_inst0 (.I(I), .O(Decode_31_8_inst0_O));
Decode_32_8 Decode_32_8_inst0 (.I(I), .O(Decode_32_8_inst0_O));
Decode_33_8 Decode_33_8_inst0 (.I(I), .O(Decode_33_8_inst0_O));
Decode_34_8 Decode_34_8_inst0 (.I(I), .O(Decode_34_8_inst0_O));
Decode_35_8 Decode_35_8_inst0 (.I(I), .O(Decode_35_8_inst0_O));
Decode_36_8 Decode_36_8_inst0 (.I(I), .O(Decode_36_8_inst0_O));
Decode_37_8 Decode_37_8_inst0 (.I(I), .O(Decode_37_8_inst0_O));
Decode_38_8 Decode_38_8_inst0 (.I(I), .O(Decode_38_8_inst0_O));
Decode_39_8 Decode_39_8_inst0 (.I(I), .O(Decode_39_8_inst0_O));
Decode_40_8 Decode_40_8_inst0 (.I(I), .O(Decode_40_8_inst0_O));
Decode_41_8 Decode_41_8_inst0 (.I(I), .O(Decode_41_8_inst0_O));
Decode_42_8 Decode_42_8_inst0 (.I(I), .O(Decode_42_8_inst0_O));
Decode_43_8 Decode_43_8_inst0 (.I(I), .O(Decode_43_8_inst0_O));
Decode_44_8 Decode_44_8_inst0 (.I(I), .O(Decode_44_8_inst0_O));
Decode_45_8 Decode_45_8_inst0 (.I(I), .O(Decode_45_8_inst0_O));
Decode_46_8 Decode_46_8_inst0 (.I(I), .O(Decode_46_8_inst0_O));
Decode_47_8 Decode_47_8_inst0 (.I(I), .O(Decode_47_8_inst0_O));
Decode_48_8 Decode_48_8_inst0 (.I(I), .O(Decode_48_8_inst0_O));
Decode_49_8 Decode_49_8_inst0 (.I(I), .O(Decode_49_8_inst0_O));
Decode_50_8 Decode_50_8_inst0 (.I(I), .O(Decode_50_8_inst0_O));
Decode_51_8 Decode_51_8_inst0 (.I(I), .O(Decode_51_8_inst0_O));
Decode_52_8 Decode_52_8_inst0 (.I(I), .O(Decode_52_8_inst0_O));
Decode_53_8 Decode_53_8_inst0 (.I(I), .O(Decode_53_8_inst0_O));
Decode_54_8 Decode_54_8_inst0 (.I(I), .O(Decode_54_8_inst0_O));
Decode_55_8 Decode_55_8_inst0 (.I(I), .O(Decode_55_8_inst0_O));
Decode_56_8 Decode_56_8_inst0 (.I(I), .O(Decode_56_8_inst0_O));
Decode_57_8 Decode_57_8_inst0 (.I(I), .O(Decode_57_8_inst0_O));
Decode_58_8 Decode_58_8_inst0 (.I(I), .O(Decode_58_8_inst0_O));
Decode_59_8 Decode_59_8_inst0 (.I(I), .O(Decode_59_8_inst0_O));
Decode_60_8 Decode_60_8_inst0 (.I(I), .O(Decode_60_8_inst0_O));
Decode_61_8 Decode_61_8_inst0 (.I(I), .O(Decode_61_8_inst0_O));
Decode_62_8 Decode_62_8_inst0 (.I(I), .O(Decode_62_8_inst0_O));
Decode_63_8 Decode_63_8_inst0 (.I(I), .O(Decode_63_8_inst0_O));
Decode_64_8 Decode_64_8_inst0 (.I(I), .O(Decode_64_8_inst0_O));
Decode_65_8 Decode_65_8_inst0 (.I(I), .O(Decode_65_8_inst0_O));
Decode_66_8 Decode_66_8_inst0 (.I(I), .O(Decode_66_8_inst0_O));
Decode_67_8 Decode_67_8_inst0 (.I(I), .O(Decode_67_8_inst0_O));
Decode_68_8 Decode_68_8_inst0 (.I(I), .O(Decode_68_8_inst0_O));
Decode_69_8 Decode_69_8_inst0 (.I(I), .O(Decode_69_8_inst0_O));
Decode_70_8 Decode_70_8_inst0 (.I(I), .O(Decode_70_8_inst0_O));
Decode_71_8 Decode_71_8_inst0 (.I(I), .O(Decode_71_8_inst0_O));
Decode_72_8 Decode_72_8_inst0 (.I(I), .O(Decode_72_8_inst0_O));
Decode_73_8 Decode_73_8_inst0 (.I(I), .O(Decode_73_8_inst0_O));
Decode_74_8 Decode_74_8_inst0 (.I(I), .O(Decode_74_8_inst0_O));
Decode_75_8 Decode_75_8_inst0 (.I(I), .O(Decode_75_8_inst0_O));
Decode_76_8 Decode_76_8_inst0 (.I(I), .O(Decode_76_8_inst0_O));
Decode_77_8 Decode_77_8_inst0 (.I(I), .O(Decode_77_8_inst0_O));
Decode_78_8 Decode_78_8_inst0 (.I(I), .O(Decode_78_8_inst0_O));
Decode_79_8 Decode_79_8_inst0 (.I(I), .O(Decode_79_8_inst0_O));
Decode_80_8 Decode_80_8_inst0 (.I(I), .O(Decode_80_8_inst0_O));
Decode_81_8 Decode_81_8_inst0 (.I(I), .O(Decode_81_8_inst0_O));
Decode_82_8 Decode_82_8_inst0 (.I(I), .O(Decode_82_8_inst0_O));
Decode_83_8 Decode_83_8_inst0 (.I(I), .O(Decode_83_8_inst0_O));
Decode_84_8 Decode_84_8_inst0 (.I(I), .O(Decode_84_8_inst0_O));
Decode_85_8 Decode_85_8_inst0 (.I(I), .O(Decode_85_8_inst0_O));
Decode_86_8 Decode_86_8_inst0 (.I(I), .O(Decode_86_8_inst0_O));
Decode_87_8 Decode_87_8_inst0 (.I(I), .O(Decode_87_8_inst0_O));
Decode_88_8 Decode_88_8_inst0 (.I(I), .O(Decode_88_8_inst0_O));
Decode_89_8 Decode_89_8_inst0 (.I(I), .O(Decode_89_8_inst0_O));
Decode_90_8 Decode_90_8_inst0 (.I(I), .O(Decode_90_8_inst0_O));
Decode_91_8 Decode_91_8_inst0 (.I(I), .O(Decode_91_8_inst0_O));
Decode_92_8 Decode_92_8_inst0 (.I(I), .O(Decode_92_8_inst0_O));
Decode_93_8 Decode_93_8_inst0 (.I(I), .O(Decode_93_8_inst0_O));
Decode_94_8 Decode_94_8_inst0 (.I(I), .O(Decode_94_8_inst0_O));
Decode_95_8 Decode_95_8_inst0 (.I(I), .O(Decode_95_8_inst0_O));
Decode_96_8 Decode_96_8_inst0 (.I(I), .O(Decode_96_8_inst0_O));
Decode_97_8 Decode_97_8_inst0 (.I(I), .O(Decode_97_8_inst0_O));
Decode_98_8 Decode_98_8_inst0 (.I(I), .O(Decode_98_8_inst0_O));
Decode_99_8 Decode_99_8_inst0 (.I(I), .O(Decode_99_8_inst0_O));
Decode_100_8 Decode_100_8_inst0 (.I(I), .O(Decode_100_8_inst0_O));
Decode_101_8 Decode_101_8_inst0 (.I(I), .O(Decode_101_8_inst0_O));
Decode_102_8 Decode_102_8_inst0 (.I(I), .O(Decode_102_8_inst0_O));
Decode_103_8 Decode_103_8_inst0 (.I(I), .O(Decode_103_8_inst0_O));
Decode_104_8 Decode_104_8_inst0 (.I(I), .O(Decode_104_8_inst0_O));
Decode_105_8 Decode_105_8_inst0 (.I(I), .O(Decode_105_8_inst0_O));
Decode_106_8 Decode_106_8_inst0 (.I(I), .O(Decode_106_8_inst0_O));
Decode_107_8 Decode_107_8_inst0 (.I(I), .O(Decode_107_8_inst0_O));
Decode_108_8 Decode_108_8_inst0 (.I(I), .O(Decode_108_8_inst0_O));
Decode_109_8 Decode_109_8_inst0 (.I(I), .O(Decode_109_8_inst0_O));
Decode_110_8 Decode_110_8_inst0 (.I(I), .O(Decode_110_8_inst0_O));
Decode_111_8 Decode_111_8_inst0 (.I(I), .O(Decode_111_8_inst0_O));
Decode_112_8 Decode_112_8_inst0 (.I(I), .O(Decode_112_8_inst0_O));
Decode_113_8 Decode_113_8_inst0 (.I(I), .O(Decode_113_8_inst0_O));
Decode_114_8 Decode_114_8_inst0 (.I(I), .O(Decode_114_8_inst0_O));
Decode_115_8 Decode_115_8_inst0 (.I(I), .O(Decode_115_8_inst0_O));
Decode_116_8 Decode_116_8_inst0 (.I(I), .O(Decode_116_8_inst0_O));
Decode_117_8 Decode_117_8_inst0 (.I(I), .O(Decode_117_8_inst0_O));
Decode_118_8 Decode_118_8_inst0 (.I(I), .O(Decode_118_8_inst0_O));
Decode_119_8 Decode_119_8_inst0 (.I(I), .O(Decode_119_8_inst0_O));
Decode_120_8 Decode_120_8_inst0 (.I(I), .O(Decode_120_8_inst0_O));
Decode_121_8 Decode_121_8_inst0 (.I(I), .O(Decode_121_8_inst0_O));
Decode_122_8 Decode_122_8_inst0 (.I(I), .O(Decode_122_8_inst0_O));
Decode_123_8 Decode_123_8_inst0 (.I(I), .O(Decode_123_8_inst0_O));
Decode_124_8 Decode_124_8_inst0 (.I(I), .O(Decode_124_8_inst0_O));
Decode_125_8 Decode_125_8_inst0 (.I(I), .O(Decode_125_8_inst0_O));
Decode_126_8 Decode_126_8_inst0 (.I(I), .O(Decode_126_8_inst0_O));
Decode_127_8 Decode_127_8_inst0 (.I(I), .O(Decode_127_8_inst0_O));
Decode_128_8 Decode_128_8_inst0 (.I(I), .O(Decode_128_8_inst0_O));
Decode_129_8 Decode_129_8_inst0 (.I(I), .O(Decode_129_8_inst0_O));
Decode_130_8 Decode_130_8_inst0 (.I(I), .O(Decode_130_8_inst0_O));
Decode_131_8 Decode_131_8_inst0 (.I(I), .O(Decode_131_8_inst0_O));
Decode_132_8 Decode_132_8_inst0 (.I(I), .O(Decode_132_8_inst0_O));
Decode_133_8 Decode_133_8_inst0 (.I(I), .O(Decode_133_8_inst0_O));
Decode_134_8 Decode_134_8_inst0 (.I(I), .O(Decode_134_8_inst0_O));
Decode_135_8 Decode_135_8_inst0 (.I(I), .O(Decode_135_8_inst0_O));
Decode_136_8 Decode_136_8_inst0 (.I(I), .O(Decode_136_8_inst0_O));
Decode_137_8 Decode_137_8_inst0 (.I(I), .O(Decode_137_8_inst0_O));
Decode_138_8 Decode_138_8_inst0 (.I(I), .O(Decode_138_8_inst0_O));
Decode_139_8 Decode_139_8_inst0 (.I(I), .O(Decode_139_8_inst0_O));
Decode_140_8 Decode_140_8_inst0 (.I(I), .O(Decode_140_8_inst0_O));
Decode_141_8 Decode_141_8_inst0 (.I(I), .O(Decode_141_8_inst0_O));
Decode_142_8 Decode_142_8_inst0 (.I(I), .O(Decode_142_8_inst0_O));
Decode_143_8 Decode_143_8_inst0 (.I(I), .O(Decode_143_8_inst0_O));
Decode_144_8 Decode_144_8_inst0 (.I(I), .O(Decode_144_8_inst0_O));
Decode_145_8 Decode_145_8_inst0 (.I(I), .O(Decode_145_8_inst0_O));
Decode_146_8 Decode_146_8_inst0 (.I(I), .O(Decode_146_8_inst0_O));
Decode_147_8 Decode_147_8_inst0 (.I(I), .O(Decode_147_8_inst0_O));
Decode_148_8 Decode_148_8_inst0 (.I(I), .O(Decode_148_8_inst0_O));
Decode_149_8 Decode_149_8_inst0 (.I(I), .O(Decode_149_8_inst0_O));
Decode_150_8 Decode_150_8_inst0 (.I(I), .O(Decode_150_8_inst0_O));
Decode_151_8 Decode_151_8_inst0 (.I(I), .O(Decode_151_8_inst0_O));
Decode_152_8 Decode_152_8_inst0 (.I(I), .O(Decode_152_8_inst0_O));
Decode_153_8 Decode_153_8_inst0 (.I(I), .O(Decode_153_8_inst0_O));
Decode_154_8 Decode_154_8_inst0 (.I(I), .O(Decode_154_8_inst0_O));
Decode_155_8 Decode_155_8_inst0 (.I(I), .O(Decode_155_8_inst0_O));
Decode_156_8 Decode_156_8_inst0 (.I(I), .O(Decode_156_8_inst0_O));
Decode_157_8 Decode_157_8_inst0 (.I(I), .O(Decode_157_8_inst0_O));
Decode_158_8 Decode_158_8_inst0 (.I(I), .O(Decode_158_8_inst0_O));
Decode_159_8 Decode_159_8_inst0 (.I(I), .O(Decode_159_8_inst0_O));
Decode_160_8 Decode_160_8_inst0 (.I(I), .O(Decode_160_8_inst0_O));
Decode_161_8 Decode_161_8_inst0 (.I(I), .O(Decode_161_8_inst0_O));
Decode_162_8 Decode_162_8_inst0 (.I(I), .O(Decode_162_8_inst0_O));
Decode_163_8 Decode_163_8_inst0 (.I(I), .O(Decode_163_8_inst0_O));
Decode_164_8 Decode_164_8_inst0 (.I(I), .O(Decode_164_8_inst0_O));
Decode_165_8 Decode_165_8_inst0 (.I(I), .O(Decode_165_8_inst0_O));
Decode_166_8 Decode_166_8_inst0 (.I(I), .O(Decode_166_8_inst0_O));
Decode_167_8 Decode_167_8_inst0 (.I(I), .O(Decode_167_8_inst0_O));
Decode_168_8 Decode_168_8_inst0 (.I(I), .O(Decode_168_8_inst0_O));
Decode_169_8 Decode_169_8_inst0 (.I(I), .O(Decode_169_8_inst0_O));
Decode_170_8 Decode_170_8_inst0 (.I(I), .O(Decode_170_8_inst0_O));
Decode_171_8 Decode_171_8_inst0 (.I(I), .O(Decode_171_8_inst0_O));
Decode_172_8 Decode_172_8_inst0 (.I(I), .O(Decode_172_8_inst0_O));
Decode_173_8 Decode_173_8_inst0 (.I(I), .O(Decode_173_8_inst0_O));
Decode_174_8 Decode_174_8_inst0 (.I(I), .O(Decode_174_8_inst0_O));
Decode_175_8 Decode_175_8_inst0 (.I(I), .O(Decode_175_8_inst0_O));
Decode_176_8 Decode_176_8_inst0 (.I(I), .O(Decode_176_8_inst0_O));
Decode_177_8 Decode_177_8_inst0 (.I(I), .O(Decode_177_8_inst0_O));
Decode_178_8 Decode_178_8_inst0 (.I(I), .O(Decode_178_8_inst0_O));
Decode_179_8 Decode_179_8_inst0 (.I(I), .O(Decode_179_8_inst0_O));
Decode_180_8 Decode_180_8_inst0 (.I(I), .O(Decode_180_8_inst0_O));
Decode_181_8 Decode_181_8_inst0 (.I(I), .O(Decode_181_8_inst0_O));
Decode_182_8 Decode_182_8_inst0 (.I(I), .O(Decode_182_8_inst0_O));
Decode_183_8 Decode_183_8_inst0 (.I(I), .O(Decode_183_8_inst0_O));
Decode_184_8 Decode_184_8_inst0 (.I(I), .O(Decode_184_8_inst0_O));
Decode_185_8 Decode_185_8_inst0 (.I(I), .O(Decode_185_8_inst0_O));
Decode_186_8 Decode_186_8_inst0 (.I(I), .O(Decode_186_8_inst0_O));
Decode_187_8 Decode_187_8_inst0 (.I(I), .O(Decode_187_8_inst0_O));
Decode_188_8 Decode_188_8_inst0 (.I(I), .O(Decode_188_8_inst0_O));
Decode_189_8 Decode_189_8_inst0 (.I(I), .O(Decode_189_8_inst0_O));
Decode_190_8 Decode_190_8_inst0 (.I(I), .O(Decode_190_8_inst0_O));
Decode_191_8 Decode_191_8_inst0 (.I(I), .O(Decode_191_8_inst0_O));
Decode_192_8 Decode_192_8_inst0 (.I(I), .O(Decode_192_8_inst0_O));
Decode_193_8 Decode_193_8_inst0 (.I(I), .O(Decode_193_8_inst0_O));
Decode_194_8 Decode_194_8_inst0 (.I(I), .O(Decode_194_8_inst0_O));
Decode_195_8 Decode_195_8_inst0 (.I(I), .O(Decode_195_8_inst0_O));
Decode_196_8 Decode_196_8_inst0 (.I(I), .O(Decode_196_8_inst0_O));
Decode_197_8 Decode_197_8_inst0 (.I(I), .O(Decode_197_8_inst0_O));
Decode_198_8 Decode_198_8_inst0 (.I(I), .O(Decode_198_8_inst0_O));
Decode_199_8 Decode_199_8_inst0 (.I(I), .O(Decode_199_8_inst0_O));
Decode_200_8 Decode_200_8_inst0 (.I(I), .O(Decode_200_8_inst0_O));
Decode_201_8 Decode_201_8_inst0 (.I(I), .O(Decode_201_8_inst0_O));
Decode_202_8 Decode_202_8_inst0 (.I(I), .O(Decode_202_8_inst0_O));
Decode_203_8 Decode_203_8_inst0 (.I(I), .O(Decode_203_8_inst0_O));
Decode_204_8 Decode_204_8_inst0 (.I(I), .O(Decode_204_8_inst0_O));
Decode_205_8 Decode_205_8_inst0 (.I(I), .O(Decode_205_8_inst0_O));
Decode_206_8 Decode_206_8_inst0 (.I(I), .O(Decode_206_8_inst0_O));
Decode_207_8 Decode_207_8_inst0 (.I(I), .O(Decode_207_8_inst0_O));
Decode_208_8 Decode_208_8_inst0 (.I(I), .O(Decode_208_8_inst0_O));
Decode_209_8 Decode_209_8_inst0 (.I(I), .O(Decode_209_8_inst0_O));
Decode_210_8 Decode_210_8_inst0 (.I(I), .O(Decode_210_8_inst0_O));
Decode_211_8 Decode_211_8_inst0 (.I(I), .O(Decode_211_8_inst0_O));
Decode_212_8 Decode_212_8_inst0 (.I(I), .O(Decode_212_8_inst0_O));
Decode_213_8 Decode_213_8_inst0 (.I(I), .O(Decode_213_8_inst0_O));
Decode_214_8 Decode_214_8_inst0 (.I(I), .O(Decode_214_8_inst0_O));
Decode_215_8 Decode_215_8_inst0 (.I(I), .O(Decode_215_8_inst0_O));
Decode_216_8 Decode_216_8_inst0 (.I(I), .O(Decode_216_8_inst0_O));
Decode_217_8 Decode_217_8_inst0 (.I(I), .O(Decode_217_8_inst0_O));
Decode_218_8 Decode_218_8_inst0 (.I(I), .O(Decode_218_8_inst0_O));
Decode_219_8 Decode_219_8_inst0 (.I(I), .O(Decode_219_8_inst0_O));
Decode_220_8 Decode_220_8_inst0 (.I(I), .O(Decode_220_8_inst0_O));
Decode_221_8 Decode_221_8_inst0 (.I(I), .O(Decode_221_8_inst0_O));
Decode_222_8 Decode_222_8_inst0 (.I(I), .O(Decode_222_8_inst0_O));
Decode_223_8 Decode_223_8_inst0 (.I(I), .O(Decode_223_8_inst0_O));
Decode_224_8 Decode_224_8_inst0 (.I(I), .O(Decode_224_8_inst0_O));
Decode_225_8 Decode_225_8_inst0 (.I(I), .O(Decode_225_8_inst0_O));
Decode_226_8 Decode_226_8_inst0 (.I(I), .O(Decode_226_8_inst0_O));
Decode_227_8 Decode_227_8_inst0 (.I(I), .O(Decode_227_8_inst0_O));
Decode_228_8 Decode_228_8_inst0 (.I(I), .O(Decode_228_8_inst0_O));
Decode_229_8 Decode_229_8_inst0 (.I(I), .O(Decode_229_8_inst0_O));
Decode_230_8 Decode_230_8_inst0 (.I(I), .O(Decode_230_8_inst0_O));
Decode_231_8 Decode_231_8_inst0 (.I(I), .O(Decode_231_8_inst0_O));
Decode_232_8 Decode_232_8_inst0 (.I(I), .O(Decode_232_8_inst0_O));
Decode_233_8 Decode_233_8_inst0 (.I(I), .O(Decode_233_8_inst0_O));
Decode_234_8 Decode_234_8_inst0 (.I(I), .O(Decode_234_8_inst0_O));
Decode_235_8 Decode_235_8_inst0 (.I(I), .O(Decode_235_8_inst0_O));
Decode_236_8 Decode_236_8_inst0 (.I(I), .O(Decode_236_8_inst0_O));
Decode_237_8 Decode_237_8_inst0 (.I(I), .O(Decode_237_8_inst0_O));
Decode_238_8 Decode_238_8_inst0 (.I(I), .O(Decode_238_8_inst0_O));
Decode_239_8 Decode_239_8_inst0 (.I(I), .O(Decode_239_8_inst0_O));
Decode_240_8 Decode_240_8_inst0 (.I(I), .O(Decode_240_8_inst0_O));
Decode_241_8 Decode_241_8_inst0 (.I(I), .O(Decode_241_8_inst0_O));
Decode_242_8 Decode_242_8_inst0 (.I(I), .O(Decode_242_8_inst0_O));
Decode_243_8 Decode_243_8_inst0 (.I(I), .O(Decode_243_8_inst0_O));
Decode_244_8 Decode_244_8_inst0 (.I(I), .O(Decode_244_8_inst0_O));
Decode_245_8 Decode_245_8_inst0 (.I(I), .O(Decode_245_8_inst0_O));
Decode_246_8 Decode_246_8_inst0 (.I(I), .O(Decode_246_8_inst0_O));
Decode_247_8 Decode_247_8_inst0 (.I(I), .O(Decode_247_8_inst0_O));
Decode_248_8 Decode_248_8_inst0 (.I(I), .O(Decode_248_8_inst0_O));
Decode_249_8 Decode_249_8_inst0 (.I(I), .O(Decode_249_8_inst0_O));
Decode_250_8 Decode_250_8_inst0 (.I(I), .O(Decode_250_8_inst0_O));
Decode_251_8 Decode_251_8_inst0 (.I(I), .O(Decode_251_8_inst0_O));
Decode_252_8 Decode_252_8_inst0 (.I(I), .O(Decode_252_8_inst0_O));
Decode_253_8 Decode_253_8_inst0 (.I(I), .O(Decode_253_8_inst0_O));
Decode_254_8 Decode_254_8_inst0 (.I(I), .O(Decode_254_8_inst0_O));
Decode_255_8 Decode_255_8_inst0 (.I(I), .O(Decode_255_8_inst0_O));
assign O = {Decode_255_8_inst0_O,Decode_254_8_inst0_O,Decode_253_8_inst0_O,Decode_252_8_inst0_O,Decode_251_8_inst0_O,Decode_250_8_inst0_O,Decode_249_8_inst0_O,Decode_248_8_inst0_O,Decode_247_8_inst0_O,Decode_246_8_inst0_O,Decode_245_8_inst0_O,Decode_244_8_inst0_O,Decode_243_8_inst0_O,Decode_242_8_inst0_O,Decode_241_8_inst0_O,Decode_240_8_inst0_O,Decode_239_8_inst0_O,Decode_238_8_inst0_O,Decode_237_8_inst0_O,Decode_236_8_inst0_O,Decode_235_8_inst0_O,Decode_234_8_inst0_O,Decode_233_8_inst0_O,Decode_232_8_inst0_O,Decode_231_8_inst0_O,Decode_230_8_inst0_O,Decode_229_8_inst0_O,Decode_228_8_inst0_O,Decode_227_8_inst0_O,Decode_226_8_inst0_O,Decode_225_8_inst0_O,Decode_224_8_inst0_O,Decode_223_8_inst0_O,Decode_222_8_inst0_O,Decode_221_8_inst0_O,Decode_220_8_inst0_O,Decode_219_8_inst0_O,Decode_218_8_inst0_O,Decode_217_8_inst0_O,Decode_216_8_inst0_O,Decode_215_8_inst0_O,Decode_214_8_inst0_O,Decode_213_8_inst0_O,Decode_212_8_inst0_O,Decode_211_8_inst0_O,Decode_210_8_inst0_O,Decode_209_8_inst0_O,Decode_208_8_inst0_O,Decode_207_8_inst0_O,Decode_206_8_inst0_O,Decode_205_8_inst0_O,Decode_204_8_inst0_O,Decode_203_8_inst0_O,Decode_202_8_inst0_O,Decode_201_8_inst0_O,Decode_200_8_inst0_O,Decode_199_8_inst0_O,Decode_198_8_inst0_O,Decode_197_8_inst0_O,Decode_196_8_inst0_O,Decode_195_8_inst0_O,Decode_194_8_inst0_O,Decode_193_8_inst0_O,Decode_192_8_inst0_O,Decode_191_8_inst0_O,Decode_190_8_inst0_O,Decode_189_8_inst0_O,Decode_188_8_inst0_O,Decode_187_8_inst0_O,Decode_186_8_inst0_O,Decode_185_8_inst0_O,Decode_184_8_inst0_O,Decode_183_8_inst0_O,Decode_182_8_inst0_O,Decode_181_8_inst0_O,Decode_180_8_inst0_O,Decode_179_8_inst0_O,Decode_178_8_inst0_O,Decode_177_8_inst0_O,Decode_176_8_inst0_O,Decode_175_8_inst0_O,Decode_174_8_inst0_O,Decode_173_8_inst0_O,Decode_172_8_inst0_O,Decode_171_8_inst0_O,Decode_170_8_inst0_O,Decode_169_8_inst0_O,Decode_168_8_inst0_O,Decode_167_8_inst0_O,Decode_166_8_inst0_O,Decode_165_8_inst0_O,Decode_164_8_inst0_O,Decode_163_8_inst0_O,Decode_162_8_inst0_O,Decode_161_8_inst0_O,Decode_160_8_inst0_O,Decode_159_8_inst0_O,Decode_158_8_inst0_O,Decode_157_8_inst0_O,Decode_156_8_inst0_O,Decode_155_8_inst0_O,Decode_154_8_inst0_O,Decode_153_8_inst0_O,Decode_152_8_inst0_O,Decode_151_8_inst0_O,Decode_150_8_inst0_O,Decode_149_8_inst0_O,Decode_148_8_inst0_O,Decode_147_8_inst0_O,Decode_146_8_inst0_O,Decode_145_8_inst0_O,Decode_144_8_inst0_O,Decode_143_8_inst0_O,Decode_142_8_inst0_O,Decode_141_8_inst0_O,Decode_140_8_inst0_O,Decode_139_8_inst0_O,Decode_138_8_inst0_O,Decode_137_8_inst0_O,Decode_136_8_inst0_O,Decode_135_8_inst0_O,Decode_134_8_inst0_O,Decode_133_8_inst0_O,Decode_132_8_inst0_O,Decode_131_8_inst0_O,Decode_130_8_inst0_O,Decode_129_8_inst0_O,Decode_128_8_inst0_O,Decode_127_8_inst0_O,Decode_126_8_inst0_O,Decode_125_8_inst0_O,Decode_124_8_inst0_O,Decode_123_8_inst0_O,Decode_122_8_inst0_O,Decode_121_8_inst0_O,Decode_120_8_inst0_O,Decode_119_8_inst0_O,Decode_118_8_inst0_O,Decode_117_8_inst0_O,Decode_116_8_inst0_O,Decode_115_8_inst0_O,Decode_114_8_inst0_O,Decode_113_8_inst0_O,Decode_112_8_inst0_O,Decode_111_8_inst0_O,Decode_110_8_inst0_O,Decode_109_8_inst0_O,Decode_108_8_inst0_O,Decode_107_8_inst0_O,Decode_106_8_inst0_O,Decode_105_8_inst0_O,Decode_104_8_inst0_O,Decode_103_8_inst0_O,Decode_102_8_inst0_O,Decode_101_8_inst0_O,Decode_100_8_inst0_O,Decode_99_8_inst0_O,Decode_98_8_inst0_O,Decode_97_8_inst0_O,Decode_96_8_inst0_O,Decode_95_8_inst0_O,Decode_94_8_inst0_O,Decode_93_8_inst0_O,Decode_92_8_inst0_O,Decode_91_8_inst0_O,Decode_90_8_inst0_O,Decode_89_8_inst0_O,Decode_88_8_inst0_O,Decode_87_8_inst0_O,Decode_86_8_inst0_O,Decode_85_8_inst0_O,Decode_84_8_inst0_O,Decode_83_8_inst0_O,Decode_82_8_inst0_O,Decode_81_8_inst0_O,Decode_80_8_inst0_O,Decode_79_8_inst0_O,Decode_78_8_inst0_O,Decode_77_8_inst0_O,Decode_76_8_inst0_O,Decode_75_8_inst0_O,Decode_74_8_inst0_O,Decode_73_8_inst0_O,Decode_72_8_inst0_O,Decode_71_8_inst0_O,Decode_70_8_inst0_O,Decode_69_8_inst0_O,Decode_68_8_inst0_O,Decode_67_8_inst0_O,Decode_66_8_inst0_O,Decode_65_8_inst0_O,Decode_64_8_inst0_O,Decode_63_8_inst0_O,Decode_62_8_inst0_O,Decode_61_8_inst0_O,Decode_60_8_inst0_O,Decode_59_8_inst0_O,Decode_58_8_inst0_O,Decode_57_8_inst0_O,Decode_56_8_inst0_O,Decode_55_8_inst0_O,Decode_54_8_inst0_O,Decode_53_8_inst0_O,Decode_52_8_inst0_O,Decode_51_8_inst0_O,Decode_50_8_inst0_O,Decode_49_8_inst0_O,Decode_48_8_inst0_O,Decode_47_8_inst0_O,Decode_46_8_inst0_O,Decode_45_8_inst0_O,Decode_44_8_inst0_O,Decode_43_8_inst0_O,Decode_42_8_inst0_O,Decode_41_8_inst0_O,Decode_40_8_inst0_O,Decode_39_8_inst0_O,Decode_38_8_inst0_O,Decode_37_8_inst0_O,Decode_36_8_inst0_O,Decode_35_8_inst0_O,Decode_34_8_inst0_O,Decode_33_8_inst0_O,Decode_32_8_inst0_O,Decode_31_8_inst0_O,Decode_30_8_inst0_O,Decode_29_8_inst0_O,Decode_28_8_inst0_O,Decode_27_8_inst0_O,Decode_26_8_inst0_O,Decode_25_8_inst0_O,Decode_24_8_inst0_O,Decode_23_8_inst0_O,Decode_22_8_inst0_O,Decode_21_8_inst0_O,Decode_20_8_inst0_O,Decode_19_8_inst0_O,Decode_18_8_inst0_O,Decode_17_8_inst0_O,Decode_16_8_inst0_O,Decode_15_8_inst0_O,Decode_14_8_inst0_O,Decode_13_8_inst0_O,Decode_12_8_inst0_O,Decode_11_8_inst0_O,Decode_10_8_inst0_O,Decode_9_8_inst0_O,Decode_8_8_inst0_O,Decode_7_8_inst0_O,Decode_6_8_inst0_O,Decode_5_8_inst0_O,Decode_4_8_inst0_O,Decode_3_8_inst0_O,Decode_2_8_inst0_O,Decode_1_8_inst0_O,Decode_0_8_inst0_O};
endmodule

