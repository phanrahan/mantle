module EQ8 (input [7:0] I0, input [7:0] I1, output  O);
wire  SB_LUT4_inst0_O;
wire  SB_LUT4_inst1_O;
wire  SB_LUT4_inst2_O;
wire  SB_LUT4_inst3_O;
wire  SB_LUT4_inst4_O;
wire  SB_LUT4_inst5_O;
wire  SB_LUT4_inst6_O;
wire  SB_LUT4_inst7_O;
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst0 (.I0(1'b1), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(SB_LUT4_inst0_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst1 (.I0(SB_LUT4_inst0_O), .I1(I0[1]), .I2(I1[1]), .I3(1'b0), .O(SB_LUT4_inst1_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst2 (.I0(SB_LUT4_inst1_O), .I1(I0[2]), .I2(I1[2]), .I3(1'b0), .O(SB_LUT4_inst2_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst3 (.I0(SB_LUT4_inst2_O), .I1(I0[3]), .I2(I1[3]), .I3(1'b0), .O(SB_LUT4_inst3_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst4 (.I0(SB_LUT4_inst3_O), .I1(I0[4]), .I2(I1[4]), .I3(1'b0), .O(SB_LUT4_inst4_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst5 (.I0(SB_LUT4_inst4_O), .I1(I0[5]), .I2(I1[5]), .I3(1'b0), .O(SB_LUT4_inst5_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst6 (.I0(SB_LUT4_inst5_O), .I1(I0[6]), .I2(I1[6]), .I3(1'b0), .O(SB_LUT4_inst6_O));
SB_LUT4 #(.LUT_INIT(16'h8282)) SB_LUT4_inst7 (.I0(SB_LUT4_inst6_O), .I1(I0[7]), .I2(I1[7]), .I3(1'b0), .O(SB_LUT4_inst7_O));
assign O = SB_LUT4_inst7_O;
endmodule

module Decode8_0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_10 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_11 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_12 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_13 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_14 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_15 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_16 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_17 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_18 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_19 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_1F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_20 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_21 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_22 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_23 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_24 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_25 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_26 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_27 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_28 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_29 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_2F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_30 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_31 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_32 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_33 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_34 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_35 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_36 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_37 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_38 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_39 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_3F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_40 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_41 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_42 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_43 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_44 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_45 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_46 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_47 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_48 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_49 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_4F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_50 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_51 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_52 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_53 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_54 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_55 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_56 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_57 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_58 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_59 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_5F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_60 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_61 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_62 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_63 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_64 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_65 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_66 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_67 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_68 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_69 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_6F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_70 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_71 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_72 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_73 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_74 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_75 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_76 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_77 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_78 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_79 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_7F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_80 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_81 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_82 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_83 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_84 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_85 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_86 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_87 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_88 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_89 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_8F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_90 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_91 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_92 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_93 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_94 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_95 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_96 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_97 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_98 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_99 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9A (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9B (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9C (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9D (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9E (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_9F (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_A9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AD (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_AF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_B9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BD (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_BF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_C9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CD (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_CF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_D9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DD (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_DF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_E9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_EA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_EB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_EC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_ED (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_EE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_EF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F0 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F1 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F2 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F3 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F4 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F5 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F6 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F7 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F8 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_F9 (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FA (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FB (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FC (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FD (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FE (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decode8_FF (input [7:0] I, output  O);
wire  EQ8_inst0_O;
EQ8 EQ8_inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(EQ8_inst0_O));
assign O = EQ8_inst0_O;
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire  Decode8_0_inst0_O;
wire  Decode8_1_inst0_O;
wire  Decode8_2_inst0_O;
wire  Decode8_3_inst0_O;
wire  Decode8_4_inst0_O;
wire  Decode8_5_inst0_O;
wire  Decode8_6_inst0_O;
wire  Decode8_7_inst0_O;
wire  Decode8_8_inst0_O;
wire  Decode8_9_inst0_O;
wire  Decode8_A_inst0_O;
wire  Decode8_B_inst0_O;
wire  Decode8_C_inst0_O;
wire  Decode8_D_inst0_O;
wire  Decode8_E_inst0_O;
wire  Decode8_F_inst0_O;
wire  Decode8_10_inst0_O;
wire  Decode8_11_inst0_O;
wire  Decode8_12_inst0_O;
wire  Decode8_13_inst0_O;
wire  Decode8_14_inst0_O;
wire  Decode8_15_inst0_O;
wire  Decode8_16_inst0_O;
wire  Decode8_17_inst0_O;
wire  Decode8_18_inst0_O;
wire  Decode8_19_inst0_O;
wire  Decode8_1A_inst0_O;
wire  Decode8_1B_inst0_O;
wire  Decode8_1C_inst0_O;
wire  Decode8_1D_inst0_O;
wire  Decode8_1E_inst0_O;
wire  Decode8_1F_inst0_O;
wire  Decode8_20_inst0_O;
wire  Decode8_21_inst0_O;
wire  Decode8_22_inst0_O;
wire  Decode8_23_inst0_O;
wire  Decode8_24_inst0_O;
wire  Decode8_25_inst0_O;
wire  Decode8_26_inst0_O;
wire  Decode8_27_inst0_O;
wire  Decode8_28_inst0_O;
wire  Decode8_29_inst0_O;
wire  Decode8_2A_inst0_O;
wire  Decode8_2B_inst0_O;
wire  Decode8_2C_inst0_O;
wire  Decode8_2D_inst0_O;
wire  Decode8_2E_inst0_O;
wire  Decode8_2F_inst0_O;
wire  Decode8_30_inst0_O;
wire  Decode8_31_inst0_O;
wire  Decode8_32_inst0_O;
wire  Decode8_33_inst0_O;
wire  Decode8_34_inst0_O;
wire  Decode8_35_inst0_O;
wire  Decode8_36_inst0_O;
wire  Decode8_37_inst0_O;
wire  Decode8_38_inst0_O;
wire  Decode8_39_inst0_O;
wire  Decode8_3A_inst0_O;
wire  Decode8_3B_inst0_O;
wire  Decode8_3C_inst0_O;
wire  Decode8_3D_inst0_O;
wire  Decode8_3E_inst0_O;
wire  Decode8_3F_inst0_O;
wire  Decode8_40_inst0_O;
wire  Decode8_41_inst0_O;
wire  Decode8_42_inst0_O;
wire  Decode8_43_inst0_O;
wire  Decode8_44_inst0_O;
wire  Decode8_45_inst0_O;
wire  Decode8_46_inst0_O;
wire  Decode8_47_inst0_O;
wire  Decode8_48_inst0_O;
wire  Decode8_49_inst0_O;
wire  Decode8_4A_inst0_O;
wire  Decode8_4B_inst0_O;
wire  Decode8_4C_inst0_O;
wire  Decode8_4D_inst0_O;
wire  Decode8_4E_inst0_O;
wire  Decode8_4F_inst0_O;
wire  Decode8_50_inst0_O;
wire  Decode8_51_inst0_O;
wire  Decode8_52_inst0_O;
wire  Decode8_53_inst0_O;
wire  Decode8_54_inst0_O;
wire  Decode8_55_inst0_O;
wire  Decode8_56_inst0_O;
wire  Decode8_57_inst0_O;
wire  Decode8_58_inst0_O;
wire  Decode8_59_inst0_O;
wire  Decode8_5A_inst0_O;
wire  Decode8_5B_inst0_O;
wire  Decode8_5C_inst0_O;
wire  Decode8_5D_inst0_O;
wire  Decode8_5E_inst0_O;
wire  Decode8_5F_inst0_O;
wire  Decode8_60_inst0_O;
wire  Decode8_61_inst0_O;
wire  Decode8_62_inst0_O;
wire  Decode8_63_inst0_O;
wire  Decode8_64_inst0_O;
wire  Decode8_65_inst0_O;
wire  Decode8_66_inst0_O;
wire  Decode8_67_inst0_O;
wire  Decode8_68_inst0_O;
wire  Decode8_69_inst0_O;
wire  Decode8_6A_inst0_O;
wire  Decode8_6B_inst0_O;
wire  Decode8_6C_inst0_O;
wire  Decode8_6D_inst0_O;
wire  Decode8_6E_inst0_O;
wire  Decode8_6F_inst0_O;
wire  Decode8_70_inst0_O;
wire  Decode8_71_inst0_O;
wire  Decode8_72_inst0_O;
wire  Decode8_73_inst0_O;
wire  Decode8_74_inst0_O;
wire  Decode8_75_inst0_O;
wire  Decode8_76_inst0_O;
wire  Decode8_77_inst0_O;
wire  Decode8_78_inst0_O;
wire  Decode8_79_inst0_O;
wire  Decode8_7A_inst0_O;
wire  Decode8_7B_inst0_O;
wire  Decode8_7C_inst0_O;
wire  Decode8_7D_inst0_O;
wire  Decode8_7E_inst0_O;
wire  Decode8_7F_inst0_O;
wire  Decode8_80_inst0_O;
wire  Decode8_81_inst0_O;
wire  Decode8_82_inst0_O;
wire  Decode8_83_inst0_O;
wire  Decode8_84_inst0_O;
wire  Decode8_85_inst0_O;
wire  Decode8_86_inst0_O;
wire  Decode8_87_inst0_O;
wire  Decode8_88_inst0_O;
wire  Decode8_89_inst0_O;
wire  Decode8_8A_inst0_O;
wire  Decode8_8B_inst0_O;
wire  Decode8_8C_inst0_O;
wire  Decode8_8D_inst0_O;
wire  Decode8_8E_inst0_O;
wire  Decode8_8F_inst0_O;
wire  Decode8_90_inst0_O;
wire  Decode8_91_inst0_O;
wire  Decode8_92_inst0_O;
wire  Decode8_93_inst0_O;
wire  Decode8_94_inst0_O;
wire  Decode8_95_inst0_O;
wire  Decode8_96_inst0_O;
wire  Decode8_97_inst0_O;
wire  Decode8_98_inst0_O;
wire  Decode8_99_inst0_O;
wire  Decode8_9A_inst0_O;
wire  Decode8_9B_inst0_O;
wire  Decode8_9C_inst0_O;
wire  Decode8_9D_inst0_O;
wire  Decode8_9E_inst0_O;
wire  Decode8_9F_inst0_O;
wire  Decode8_A0_inst0_O;
wire  Decode8_A1_inst0_O;
wire  Decode8_A2_inst0_O;
wire  Decode8_A3_inst0_O;
wire  Decode8_A4_inst0_O;
wire  Decode8_A5_inst0_O;
wire  Decode8_A6_inst0_O;
wire  Decode8_A7_inst0_O;
wire  Decode8_A8_inst0_O;
wire  Decode8_A9_inst0_O;
wire  Decode8_AA_inst0_O;
wire  Decode8_AB_inst0_O;
wire  Decode8_AC_inst0_O;
wire  Decode8_AD_inst0_O;
wire  Decode8_AE_inst0_O;
wire  Decode8_AF_inst0_O;
wire  Decode8_B0_inst0_O;
wire  Decode8_B1_inst0_O;
wire  Decode8_B2_inst0_O;
wire  Decode8_B3_inst0_O;
wire  Decode8_B4_inst0_O;
wire  Decode8_B5_inst0_O;
wire  Decode8_B6_inst0_O;
wire  Decode8_B7_inst0_O;
wire  Decode8_B8_inst0_O;
wire  Decode8_B9_inst0_O;
wire  Decode8_BA_inst0_O;
wire  Decode8_BB_inst0_O;
wire  Decode8_BC_inst0_O;
wire  Decode8_BD_inst0_O;
wire  Decode8_BE_inst0_O;
wire  Decode8_BF_inst0_O;
wire  Decode8_C0_inst0_O;
wire  Decode8_C1_inst0_O;
wire  Decode8_C2_inst0_O;
wire  Decode8_C3_inst0_O;
wire  Decode8_C4_inst0_O;
wire  Decode8_C5_inst0_O;
wire  Decode8_C6_inst0_O;
wire  Decode8_C7_inst0_O;
wire  Decode8_C8_inst0_O;
wire  Decode8_C9_inst0_O;
wire  Decode8_CA_inst0_O;
wire  Decode8_CB_inst0_O;
wire  Decode8_CC_inst0_O;
wire  Decode8_CD_inst0_O;
wire  Decode8_CE_inst0_O;
wire  Decode8_CF_inst0_O;
wire  Decode8_D0_inst0_O;
wire  Decode8_D1_inst0_O;
wire  Decode8_D2_inst0_O;
wire  Decode8_D3_inst0_O;
wire  Decode8_D4_inst0_O;
wire  Decode8_D5_inst0_O;
wire  Decode8_D6_inst0_O;
wire  Decode8_D7_inst0_O;
wire  Decode8_D8_inst0_O;
wire  Decode8_D9_inst0_O;
wire  Decode8_DA_inst0_O;
wire  Decode8_DB_inst0_O;
wire  Decode8_DC_inst0_O;
wire  Decode8_DD_inst0_O;
wire  Decode8_DE_inst0_O;
wire  Decode8_DF_inst0_O;
wire  Decode8_E0_inst0_O;
wire  Decode8_E1_inst0_O;
wire  Decode8_E2_inst0_O;
wire  Decode8_E3_inst0_O;
wire  Decode8_E4_inst0_O;
wire  Decode8_E5_inst0_O;
wire  Decode8_E6_inst0_O;
wire  Decode8_E7_inst0_O;
wire  Decode8_E8_inst0_O;
wire  Decode8_E9_inst0_O;
wire  Decode8_EA_inst0_O;
wire  Decode8_EB_inst0_O;
wire  Decode8_EC_inst0_O;
wire  Decode8_ED_inst0_O;
wire  Decode8_EE_inst0_O;
wire  Decode8_EF_inst0_O;
wire  Decode8_F0_inst0_O;
wire  Decode8_F1_inst0_O;
wire  Decode8_F2_inst0_O;
wire  Decode8_F3_inst0_O;
wire  Decode8_F4_inst0_O;
wire  Decode8_F5_inst0_O;
wire  Decode8_F6_inst0_O;
wire  Decode8_F7_inst0_O;
wire  Decode8_F8_inst0_O;
wire  Decode8_F9_inst0_O;
wire  Decode8_FA_inst0_O;
wire  Decode8_FB_inst0_O;
wire  Decode8_FC_inst0_O;
wire  Decode8_FD_inst0_O;
wire  Decode8_FE_inst0_O;
wire  Decode8_FF_inst0_O;
Decode8_0 Decode8_0_inst0 (.I(I), .O(Decode8_0_inst0_O));
Decode8_1 Decode8_1_inst0 (.I(I), .O(Decode8_1_inst0_O));
Decode8_2 Decode8_2_inst0 (.I(I), .O(Decode8_2_inst0_O));
Decode8_3 Decode8_3_inst0 (.I(I), .O(Decode8_3_inst0_O));
Decode8_4 Decode8_4_inst0 (.I(I), .O(Decode8_4_inst0_O));
Decode8_5 Decode8_5_inst0 (.I(I), .O(Decode8_5_inst0_O));
Decode8_6 Decode8_6_inst0 (.I(I), .O(Decode8_6_inst0_O));
Decode8_7 Decode8_7_inst0 (.I(I), .O(Decode8_7_inst0_O));
Decode8_8 Decode8_8_inst0 (.I(I), .O(Decode8_8_inst0_O));
Decode8_9 Decode8_9_inst0 (.I(I), .O(Decode8_9_inst0_O));
Decode8_A Decode8_A_inst0 (.I(I), .O(Decode8_A_inst0_O));
Decode8_B Decode8_B_inst0 (.I(I), .O(Decode8_B_inst0_O));
Decode8_C Decode8_C_inst0 (.I(I), .O(Decode8_C_inst0_O));
Decode8_D Decode8_D_inst0 (.I(I), .O(Decode8_D_inst0_O));
Decode8_E Decode8_E_inst0 (.I(I), .O(Decode8_E_inst0_O));
Decode8_F Decode8_F_inst0 (.I(I), .O(Decode8_F_inst0_O));
Decode8_10 Decode8_10_inst0 (.I(I), .O(Decode8_10_inst0_O));
Decode8_11 Decode8_11_inst0 (.I(I), .O(Decode8_11_inst0_O));
Decode8_12 Decode8_12_inst0 (.I(I), .O(Decode8_12_inst0_O));
Decode8_13 Decode8_13_inst0 (.I(I), .O(Decode8_13_inst0_O));
Decode8_14 Decode8_14_inst0 (.I(I), .O(Decode8_14_inst0_O));
Decode8_15 Decode8_15_inst0 (.I(I), .O(Decode8_15_inst0_O));
Decode8_16 Decode8_16_inst0 (.I(I), .O(Decode8_16_inst0_O));
Decode8_17 Decode8_17_inst0 (.I(I), .O(Decode8_17_inst0_O));
Decode8_18 Decode8_18_inst0 (.I(I), .O(Decode8_18_inst0_O));
Decode8_19 Decode8_19_inst0 (.I(I), .O(Decode8_19_inst0_O));
Decode8_1A Decode8_1A_inst0 (.I(I), .O(Decode8_1A_inst0_O));
Decode8_1B Decode8_1B_inst0 (.I(I), .O(Decode8_1B_inst0_O));
Decode8_1C Decode8_1C_inst0 (.I(I), .O(Decode8_1C_inst0_O));
Decode8_1D Decode8_1D_inst0 (.I(I), .O(Decode8_1D_inst0_O));
Decode8_1E Decode8_1E_inst0 (.I(I), .O(Decode8_1E_inst0_O));
Decode8_1F Decode8_1F_inst0 (.I(I), .O(Decode8_1F_inst0_O));
Decode8_20 Decode8_20_inst0 (.I(I), .O(Decode8_20_inst0_O));
Decode8_21 Decode8_21_inst0 (.I(I), .O(Decode8_21_inst0_O));
Decode8_22 Decode8_22_inst0 (.I(I), .O(Decode8_22_inst0_O));
Decode8_23 Decode8_23_inst0 (.I(I), .O(Decode8_23_inst0_O));
Decode8_24 Decode8_24_inst0 (.I(I), .O(Decode8_24_inst0_O));
Decode8_25 Decode8_25_inst0 (.I(I), .O(Decode8_25_inst0_O));
Decode8_26 Decode8_26_inst0 (.I(I), .O(Decode8_26_inst0_O));
Decode8_27 Decode8_27_inst0 (.I(I), .O(Decode8_27_inst0_O));
Decode8_28 Decode8_28_inst0 (.I(I), .O(Decode8_28_inst0_O));
Decode8_29 Decode8_29_inst0 (.I(I), .O(Decode8_29_inst0_O));
Decode8_2A Decode8_2A_inst0 (.I(I), .O(Decode8_2A_inst0_O));
Decode8_2B Decode8_2B_inst0 (.I(I), .O(Decode8_2B_inst0_O));
Decode8_2C Decode8_2C_inst0 (.I(I), .O(Decode8_2C_inst0_O));
Decode8_2D Decode8_2D_inst0 (.I(I), .O(Decode8_2D_inst0_O));
Decode8_2E Decode8_2E_inst0 (.I(I), .O(Decode8_2E_inst0_O));
Decode8_2F Decode8_2F_inst0 (.I(I), .O(Decode8_2F_inst0_O));
Decode8_30 Decode8_30_inst0 (.I(I), .O(Decode8_30_inst0_O));
Decode8_31 Decode8_31_inst0 (.I(I), .O(Decode8_31_inst0_O));
Decode8_32 Decode8_32_inst0 (.I(I), .O(Decode8_32_inst0_O));
Decode8_33 Decode8_33_inst0 (.I(I), .O(Decode8_33_inst0_O));
Decode8_34 Decode8_34_inst0 (.I(I), .O(Decode8_34_inst0_O));
Decode8_35 Decode8_35_inst0 (.I(I), .O(Decode8_35_inst0_O));
Decode8_36 Decode8_36_inst0 (.I(I), .O(Decode8_36_inst0_O));
Decode8_37 Decode8_37_inst0 (.I(I), .O(Decode8_37_inst0_O));
Decode8_38 Decode8_38_inst0 (.I(I), .O(Decode8_38_inst0_O));
Decode8_39 Decode8_39_inst0 (.I(I), .O(Decode8_39_inst0_O));
Decode8_3A Decode8_3A_inst0 (.I(I), .O(Decode8_3A_inst0_O));
Decode8_3B Decode8_3B_inst0 (.I(I), .O(Decode8_3B_inst0_O));
Decode8_3C Decode8_3C_inst0 (.I(I), .O(Decode8_3C_inst0_O));
Decode8_3D Decode8_3D_inst0 (.I(I), .O(Decode8_3D_inst0_O));
Decode8_3E Decode8_3E_inst0 (.I(I), .O(Decode8_3E_inst0_O));
Decode8_3F Decode8_3F_inst0 (.I(I), .O(Decode8_3F_inst0_O));
Decode8_40 Decode8_40_inst0 (.I(I), .O(Decode8_40_inst0_O));
Decode8_41 Decode8_41_inst0 (.I(I), .O(Decode8_41_inst0_O));
Decode8_42 Decode8_42_inst0 (.I(I), .O(Decode8_42_inst0_O));
Decode8_43 Decode8_43_inst0 (.I(I), .O(Decode8_43_inst0_O));
Decode8_44 Decode8_44_inst0 (.I(I), .O(Decode8_44_inst0_O));
Decode8_45 Decode8_45_inst0 (.I(I), .O(Decode8_45_inst0_O));
Decode8_46 Decode8_46_inst0 (.I(I), .O(Decode8_46_inst0_O));
Decode8_47 Decode8_47_inst0 (.I(I), .O(Decode8_47_inst0_O));
Decode8_48 Decode8_48_inst0 (.I(I), .O(Decode8_48_inst0_O));
Decode8_49 Decode8_49_inst0 (.I(I), .O(Decode8_49_inst0_O));
Decode8_4A Decode8_4A_inst0 (.I(I), .O(Decode8_4A_inst0_O));
Decode8_4B Decode8_4B_inst0 (.I(I), .O(Decode8_4B_inst0_O));
Decode8_4C Decode8_4C_inst0 (.I(I), .O(Decode8_4C_inst0_O));
Decode8_4D Decode8_4D_inst0 (.I(I), .O(Decode8_4D_inst0_O));
Decode8_4E Decode8_4E_inst0 (.I(I), .O(Decode8_4E_inst0_O));
Decode8_4F Decode8_4F_inst0 (.I(I), .O(Decode8_4F_inst0_O));
Decode8_50 Decode8_50_inst0 (.I(I), .O(Decode8_50_inst0_O));
Decode8_51 Decode8_51_inst0 (.I(I), .O(Decode8_51_inst0_O));
Decode8_52 Decode8_52_inst0 (.I(I), .O(Decode8_52_inst0_O));
Decode8_53 Decode8_53_inst0 (.I(I), .O(Decode8_53_inst0_O));
Decode8_54 Decode8_54_inst0 (.I(I), .O(Decode8_54_inst0_O));
Decode8_55 Decode8_55_inst0 (.I(I), .O(Decode8_55_inst0_O));
Decode8_56 Decode8_56_inst0 (.I(I), .O(Decode8_56_inst0_O));
Decode8_57 Decode8_57_inst0 (.I(I), .O(Decode8_57_inst0_O));
Decode8_58 Decode8_58_inst0 (.I(I), .O(Decode8_58_inst0_O));
Decode8_59 Decode8_59_inst0 (.I(I), .O(Decode8_59_inst0_O));
Decode8_5A Decode8_5A_inst0 (.I(I), .O(Decode8_5A_inst0_O));
Decode8_5B Decode8_5B_inst0 (.I(I), .O(Decode8_5B_inst0_O));
Decode8_5C Decode8_5C_inst0 (.I(I), .O(Decode8_5C_inst0_O));
Decode8_5D Decode8_5D_inst0 (.I(I), .O(Decode8_5D_inst0_O));
Decode8_5E Decode8_5E_inst0 (.I(I), .O(Decode8_5E_inst0_O));
Decode8_5F Decode8_5F_inst0 (.I(I), .O(Decode8_5F_inst0_O));
Decode8_60 Decode8_60_inst0 (.I(I), .O(Decode8_60_inst0_O));
Decode8_61 Decode8_61_inst0 (.I(I), .O(Decode8_61_inst0_O));
Decode8_62 Decode8_62_inst0 (.I(I), .O(Decode8_62_inst0_O));
Decode8_63 Decode8_63_inst0 (.I(I), .O(Decode8_63_inst0_O));
Decode8_64 Decode8_64_inst0 (.I(I), .O(Decode8_64_inst0_O));
Decode8_65 Decode8_65_inst0 (.I(I), .O(Decode8_65_inst0_O));
Decode8_66 Decode8_66_inst0 (.I(I), .O(Decode8_66_inst0_O));
Decode8_67 Decode8_67_inst0 (.I(I), .O(Decode8_67_inst0_O));
Decode8_68 Decode8_68_inst0 (.I(I), .O(Decode8_68_inst0_O));
Decode8_69 Decode8_69_inst0 (.I(I), .O(Decode8_69_inst0_O));
Decode8_6A Decode8_6A_inst0 (.I(I), .O(Decode8_6A_inst0_O));
Decode8_6B Decode8_6B_inst0 (.I(I), .O(Decode8_6B_inst0_O));
Decode8_6C Decode8_6C_inst0 (.I(I), .O(Decode8_6C_inst0_O));
Decode8_6D Decode8_6D_inst0 (.I(I), .O(Decode8_6D_inst0_O));
Decode8_6E Decode8_6E_inst0 (.I(I), .O(Decode8_6E_inst0_O));
Decode8_6F Decode8_6F_inst0 (.I(I), .O(Decode8_6F_inst0_O));
Decode8_70 Decode8_70_inst0 (.I(I), .O(Decode8_70_inst0_O));
Decode8_71 Decode8_71_inst0 (.I(I), .O(Decode8_71_inst0_O));
Decode8_72 Decode8_72_inst0 (.I(I), .O(Decode8_72_inst0_O));
Decode8_73 Decode8_73_inst0 (.I(I), .O(Decode8_73_inst0_O));
Decode8_74 Decode8_74_inst0 (.I(I), .O(Decode8_74_inst0_O));
Decode8_75 Decode8_75_inst0 (.I(I), .O(Decode8_75_inst0_O));
Decode8_76 Decode8_76_inst0 (.I(I), .O(Decode8_76_inst0_O));
Decode8_77 Decode8_77_inst0 (.I(I), .O(Decode8_77_inst0_O));
Decode8_78 Decode8_78_inst0 (.I(I), .O(Decode8_78_inst0_O));
Decode8_79 Decode8_79_inst0 (.I(I), .O(Decode8_79_inst0_O));
Decode8_7A Decode8_7A_inst0 (.I(I), .O(Decode8_7A_inst0_O));
Decode8_7B Decode8_7B_inst0 (.I(I), .O(Decode8_7B_inst0_O));
Decode8_7C Decode8_7C_inst0 (.I(I), .O(Decode8_7C_inst0_O));
Decode8_7D Decode8_7D_inst0 (.I(I), .O(Decode8_7D_inst0_O));
Decode8_7E Decode8_7E_inst0 (.I(I), .O(Decode8_7E_inst0_O));
Decode8_7F Decode8_7F_inst0 (.I(I), .O(Decode8_7F_inst0_O));
Decode8_80 Decode8_80_inst0 (.I(I), .O(Decode8_80_inst0_O));
Decode8_81 Decode8_81_inst0 (.I(I), .O(Decode8_81_inst0_O));
Decode8_82 Decode8_82_inst0 (.I(I), .O(Decode8_82_inst0_O));
Decode8_83 Decode8_83_inst0 (.I(I), .O(Decode8_83_inst0_O));
Decode8_84 Decode8_84_inst0 (.I(I), .O(Decode8_84_inst0_O));
Decode8_85 Decode8_85_inst0 (.I(I), .O(Decode8_85_inst0_O));
Decode8_86 Decode8_86_inst0 (.I(I), .O(Decode8_86_inst0_O));
Decode8_87 Decode8_87_inst0 (.I(I), .O(Decode8_87_inst0_O));
Decode8_88 Decode8_88_inst0 (.I(I), .O(Decode8_88_inst0_O));
Decode8_89 Decode8_89_inst0 (.I(I), .O(Decode8_89_inst0_O));
Decode8_8A Decode8_8A_inst0 (.I(I), .O(Decode8_8A_inst0_O));
Decode8_8B Decode8_8B_inst0 (.I(I), .O(Decode8_8B_inst0_O));
Decode8_8C Decode8_8C_inst0 (.I(I), .O(Decode8_8C_inst0_O));
Decode8_8D Decode8_8D_inst0 (.I(I), .O(Decode8_8D_inst0_O));
Decode8_8E Decode8_8E_inst0 (.I(I), .O(Decode8_8E_inst0_O));
Decode8_8F Decode8_8F_inst0 (.I(I), .O(Decode8_8F_inst0_O));
Decode8_90 Decode8_90_inst0 (.I(I), .O(Decode8_90_inst0_O));
Decode8_91 Decode8_91_inst0 (.I(I), .O(Decode8_91_inst0_O));
Decode8_92 Decode8_92_inst0 (.I(I), .O(Decode8_92_inst0_O));
Decode8_93 Decode8_93_inst0 (.I(I), .O(Decode8_93_inst0_O));
Decode8_94 Decode8_94_inst0 (.I(I), .O(Decode8_94_inst0_O));
Decode8_95 Decode8_95_inst0 (.I(I), .O(Decode8_95_inst0_O));
Decode8_96 Decode8_96_inst0 (.I(I), .O(Decode8_96_inst0_O));
Decode8_97 Decode8_97_inst0 (.I(I), .O(Decode8_97_inst0_O));
Decode8_98 Decode8_98_inst0 (.I(I), .O(Decode8_98_inst0_O));
Decode8_99 Decode8_99_inst0 (.I(I), .O(Decode8_99_inst0_O));
Decode8_9A Decode8_9A_inst0 (.I(I), .O(Decode8_9A_inst0_O));
Decode8_9B Decode8_9B_inst0 (.I(I), .O(Decode8_9B_inst0_O));
Decode8_9C Decode8_9C_inst0 (.I(I), .O(Decode8_9C_inst0_O));
Decode8_9D Decode8_9D_inst0 (.I(I), .O(Decode8_9D_inst0_O));
Decode8_9E Decode8_9E_inst0 (.I(I), .O(Decode8_9E_inst0_O));
Decode8_9F Decode8_9F_inst0 (.I(I), .O(Decode8_9F_inst0_O));
Decode8_A0 Decode8_A0_inst0 (.I(I), .O(Decode8_A0_inst0_O));
Decode8_A1 Decode8_A1_inst0 (.I(I), .O(Decode8_A1_inst0_O));
Decode8_A2 Decode8_A2_inst0 (.I(I), .O(Decode8_A2_inst0_O));
Decode8_A3 Decode8_A3_inst0 (.I(I), .O(Decode8_A3_inst0_O));
Decode8_A4 Decode8_A4_inst0 (.I(I), .O(Decode8_A4_inst0_O));
Decode8_A5 Decode8_A5_inst0 (.I(I), .O(Decode8_A5_inst0_O));
Decode8_A6 Decode8_A6_inst0 (.I(I), .O(Decode8_A6_inst0_O));
Decode8_A7 Decode8_A7_inst0 (.I(I), .O(Decode8_A7_inst0_O));
Decode8_A8 Decode8_A8_inst0 (.I(I), .O(Decode8_A8_inst0_O));
Decode8_A9 Decode8_A9_inst0 (.I(I), .O(Decode8_A9_inst0_O));
Decode8_AA Decode8_AA_inst0 (.I(I), .O(Decode8_AA_inst0_O));
Decode8_AB Decode8_AB_inst0 (.I(I), .O(Decode8_AB_inst0_O));
Decode8_AC Decode8_AC_inst0 (.I(I), .O(Decode8_AC_inst0_O));
Decode8_AD Decode8_AD_inst0 (.I(I), .O(Decode8_AD_inst0_O));
Decode8_AE Decode8_AE_inst0 (.I(I), .O(Decode8_AE_inst0_O));
Decode8_AF Decode8_AF_inst0 (.I(I), .O(Decode8_AF_inst0_O));
Decode8_B0 Decode8_B0_inst0 (.I(I), .O(Decode8_B0_inst0_O));
Decode8_B1 Decode8_B1_inst0 (.I(I), .O(Decode8_B1_inst0_O));
Decode8_B2 Decode8_B2_inst0 (.I(I), .O(Decode8_B2_inst0_O));
Decode8_B3 Decode8_B3_inst0 (.I(I), .O(Decode8_B3_inst0_O));
Decode8_B4 Decode8_B4_inst0 (.I(I), .O(Decode8_B4_inst0_O));
Decode8_B5 Decode8_B5_inst0 (.I(I), .O(Decode8_B5_inst0_O));
Decode8_B6 Decode8_B6_inst0 (.I(I), .O(Decode8_B6_inst0_O));
Decode8_B7 Decode8_B7_inst0 (.I(I), .O(Decode8_B7_inst0_O));
Decode8_B8 Decode8_B8_inst0 (.I(I), .O(Decode8_B8_inst0_O));
Decode8_B9 Decode8_B9_inst0 (.I(I), .O(Decode8_B9_inst0_O));
Decode8_BA Decode8_BA_inst0 (.I(I), .O(Decode8_BA_inst0_O));
Decode8_BB Decode8_BB_inst0 (.I(I), .O(Decode8_BB_inst0_O));
Decode8_BC Decode8_BC_inst0 (.I(I), .O(Decode8_BC_inst0_O));
Decode8_BD Decode8_BD_inst0 (.I(I), .O(Decode8_BD_inst0_O));
Decode8_BE Decode8_BE_inst0 (.I(I), .O(Decode8_BE_inst0_O));
Decode8_BF Decode8_BF_inst0 (.I(I), .O(Decode8_BF_inst0_O));
Decode8_C0 Decode8_C0_inst0 (.I(I), .O(Decode8_C0_inst0_O));
Decode8_C1 Decode8_C1_inst0 (.I(I), .O(Decode8_C1_inst0_O));
Decode8_C2 Decode8_C2_inst0 (.I(I), .O(Decode8_C2_inst0_O));
Decode8_C3 Decode8_C3_inst0 (.I(I), .O(Decode8_C3_inst0_O));
Decode8_C4 Decode8_C4_inst0 (.I(I), .O(Decode8_C4_inst0_O));
Decode8_C5 Decode8_C5_inst0 (.I(I), .O(Decode8_C5_inst0_O));
Decode8_C6 Decode8_C6_inst0 (.I(I), .O(Decode8_C6_inst0_O));
Decode8_C7 Decode8_C7_inst0 (.I(I), .O(Decode8_C7_inst0_O));
Decode8_C8 Decode8_C8_inst0 (.I(I), .O(Decode8_C8_inst0_O));
Decode8_C9 Decode8_C9_inst0 (.I(I), .O(Decode8_C9_inst0_O));
Decode8_CA Decode8_CA_inst0 (.I(I), .O(Decode8_CA_inst0_O));
Decode8_CB Decode8_CB_inst0 (.I(I), .O(Decode8_CB_inst0_O));
Decode8_CC Decode8_CC_inst0 (.I(I), .O(Decode8_CC_inst0_O));
Decode8_CD Decode8_CD_inst0 (.I(I), .O(Decode8_CD_inst0_O));
Decode8_CE Decode8_CE_inst0 (.I(I), .O(Decode8_CE_inst0_O));
Decode8_CF Decode8_CF_inst0 (.I(I), .O(Decode8_CF_inst0_O));
Decode8_D0 Decode8_D0_inst0 (.I(I), .O(Decode8_D0_inst0_O));
Decode8_D1 Decode8_D1_inst0 (.I(I), .O(Decode8_D1_inst0_O));
Decode8_D2 Decode8_D2_inst0 (.I(I), .O(Decode8_D2_inst0_O));
Decode8_D3 Decode8_D3_inst0 (.I(I), .O(Decode8_D3_inst0_O));
Decode8_D4 Decode8_D4_inst0 (.I(I), .O(Decode8_D4_inst0_O));
Decode8_D5 Decode8_D5_inst0 (.I(I), .O(Decode8_D5_inst0_O));
Decode8_D6 Decode8_D6_inst0 (.I(I), .O(Decode8_D6_inst0_O));
Decode8_D7 Decode8_D7_inst0 (.I(I), .O(Decode8_D7_inst0_O));
Decode8_D8 Decode8_D8_inst0 (.I(I), .O(Decode8_D8_inst0_O));
Decode8_D9 Decode8_D9_inst0 (.I(I), .O(Decode8_D9_inst0_O));
Decode8_DA Decode8_DA_inst0 (.I(I), .O(Decode8_DA_inst0_O));
Decode8_DB Decode8_DB_inst0 (.I(I), .O(Decode8_DB_inst0_O));
Decode8_DC Decode8_DC_inst0 (.I(I), .O(Decode8_DC_inst0_O));
Decode8_DD Decode8_DD_inst0 (.I(I), .O(Decode8_DD_inst0_O));
Decode8_DE Decode8_DE_inst0 (.I(I), .O(Decode8_DE_inst0_O));
Decode8_DF Decode8_DF_inst0 (.I(I), .O(Decode8_DF_inst0_O));
Decode8_E0 Decode8_E0_inst0 (.I(I), .O(Decode8_E0_inst0_O));
Decode8_E1 Decode8_E1_inst0 (.I(I), .O(Decode8_E1_inst0_O));
Decode8_E2 Decode8_E2_inst0 (.I(I), .O(Decode8_E2_inst0_O));
Decode8_E3 Decode8_E3_inst0 (.I(I), .O(Decode8_E3_inst0_O));
Decode8_E4 Decode8_E4_inst0 (.I(I), .O(Decode8_E4_inst0_O));
Decode8_E5 Decode8_E5_inst0 (.I(I), .O(Decode8_E5_inst0_O));
Decode8_E6 Decode8_E6_inst0 (.I(I), .O(Decode8_E6_inst0_O));
Decode8_E7 Decode8_E7_inst0 (.I(I), .O(Decode8_E7_inst0_O));
Decode8_E8 Decode8_E8_inst0 (.I(I), .O(Decode8_E8_inst0_O));
Decode8_E9 Decode8_E9_inst0 (.I(I), .O(Decode8_E9_inst0_O));
Decode8_EA Decode8_EA_inst0 (.I(I), .O(Decode8_EA_inst0_O));
Decode8_EB Decode8_EB_inst0 (.I(I), .O(Decode8_EB_inst0_O));
Decode8_EC Decode8_EC_inst0 (.I(I), .O(Decode8_EC_inst0_O));
Decode8_ED Decode8_ED_inst0 (.I(I), .O(Decode8_ED_inst0_O));
Decode8_EE Decode8_EE_inst0 (.I(I), .O(Decode8_EE_inst0_O));
Decode8_EF Decode8_EF_inst0 (.I(I), .O(Decode8_EF_inst0_O));
Decode8_F0 Decode8_F0_inst0 (.I(I), .O(Decode8_F0_inst0_O));
Decode8_F1 Decode8_F1_inst0 (.I(I), .O(Decode8_F1_inst0_O));
Decode8_F2 Decode8_F2_inst0 (.I(I), .O(Decode8_F2_inst0_O));
Decode8_F3 Decode8_F3_inst0 (.I(I), .O(Decode8_F3_inst0_O));
Decode8_F4 Decode8_F4_inst0 (.I(I), .O(Decode8_F4_inst0_O));
Decode8_F5 Decode8_F5_inst0 (.I(I), .O(Decode8_F5_inst0_O));
Decode8_F6 Decode8_F6_inst0 (.I(I), .O(Decode8_F6_inst0_O));
Decode8_F7 Decode8_F7_inst0 (.I(I), .O(Decode8_F7_inst0_O));
Decode8_F8 Decode8_F8_inst0 (.I(I), .O(Decode8_F8_inst0_O));
Decode8_F9 Decode8_F9_inst0 (.I(I), .O(Decode8_F9_inst0_O));
Decode8_FA Decode8_FA_inst0 (.I(I), .O(Decode8_FA_inst0_O));
Decode8_FB Decode8_FB_inst0 (.I(I), .O(Decode8_FB_inst0_O));
Decode8_FC Decode8_FC_inst0 (.I(I), .O(Decode8_FC_inst0_O));
Decode8_FD Decode8_FD_inst0 (.I(I), .O(Decode8_FD_inst0_O));
Decode8_FE Decode8_FE_inst0 (.I(I), .O(Decode8_FE_inst0_O));
Decode8_FF Decode8_FF_inst0 (.I(I), .O(Decode8_FF_inst0_O));
assign O = {Decode8_FF_inst0_O,Decode8_FE_inst0_O,Decode8_FD_inst0_O,Decode8_FC_inst0_O,Decode8_FB_inst0_O,Decode8_FA_inst0_O,Decode8_F9_inst0_O,Decode8_F8_inst0_O,Decode8_F7_inst0_O,Decode8_F6_inst0_O,Decode8_F5_inst0_O,Decode8_F4_inst0_O,Decode8_F3_inst0_O,Decode8_F2_inst0_O,Decode8_F1_inst0_O,Decode8_F0_inst0_O,Decode8_EF_inst0_O,Decode8_EE_inst0_O,Decode8_ED_inst0_O,Decode8_EC_inst0_O,Decode8_EB_inst0_O,Decode8_EA_inst0_O,Decode8_E9_inst0_O,Decode8_E8_inst0_O,Decode8_E7_inst0_O,Decode8_E6_inst0_O,Decode8_E5_inst0_O,Decode8_E4_inst0_O,Decode8_E3_inst0_O,Decode8_E2_inst0_O,Decode8_E1_inst0_O,Decode8_E0_inst0_O,Decode8_DF_inst0_O,Decode8_DE_inst0_O,Decode8_DD_inst0_O,Decode8_DC_inst0_O,Decode8_DB_inst0_O,Decode8_DA_inst0_O,Decode8_D9_inst0_O,Decode8_D8_inst0_O,Decode8_D7_inst0_O,Decode8_D6_inst0_O,Decode8_D5_inst0_O,Decode8_D4_inst0_O,Decode8_D3_inst0_O,Decode8_D2_inst0_O,Decode8_D1_inst0_O,Decode8_D0_inst0_O,Decode8_CF_inst0_O,Decode8_CE_inst0_O,Decode8_CD_inst0_O,Decode8_CC_inst0_O,Decode8_CB_inst0_O,Decode8_CA_inst0_O,Decode8_C9_inst0_O,Decode8_C8_inst0_O,Decode8_C7_inst0_O,Decode8_C6_inst0_O,Decode8_C5_inst0_O,Decode8_C4_inst0_O,Decode8_C3_inst0_O,Decode8_C2_inst0_O,Decode8_C1_inst0_O,Decode8_C0_inst0_O,Decode8_BF_inst0_O,Decode8_BE_inst0_O,Decode8_BD_inst0_O,Decode8_BC_inst0_O,Decode8_BB_inst0_O,Decode8_BA_inst0_O,Decode8_B9_inst0_O,Decode8_B8_inst0_O,Decode8_B7_inst0_O,Decode8_B6_inst0_O,Decode8_B5_inst0_O,Decode8_B4_inst0_O,Decode8_B3_inst0_O,Decode8_B2_inst0_O,Decode8_B1_inst0_O,Decode8_B0_inst0_O,Decode8_AF_inst0_O,Decode8_AE_inst0_O,Decode8_AD_inst0_O,Decode8_AC_inst0_O,Decode8_AB_inst0_O,Decode8_AA_inst0_O,Decode8_A9_inst0_O,Decode8_A8_inst0_O,Decode8_A7_inst0_O,Decode8_A6_inst0_O,Decode8_A5_inst0_O,Decode8_A4_inst0_O,Decode8_A3_inst0_O,Decode8_A2_inst0_O,Decode8_A1_inst0_O,Decode8_A0_inst0_O,Decode8_9F_inst0_O,Decode8_9E_inst0_O,Decode8_9D_inst0_O,Decode8_9C_inst0_O,Decode8_9B_inst0_O,Decode8_9A_inst0_O,Decode8_99_inst0_O,Decode8_98_inst0_O,Decode8_97_inst0_O,Decode8_96_inst0_O,Decode8_95_inst0_O,Decode8_94_inst0_O,Decode8_93_inst0_O,Decode8_92_inst0_O,Decode8_91_inst0_O,Decode8_90_inst0_O,Decode8_8F_inst0_O,Decode8_8E_inst0_O,Decode8_8D_inst0_O,Decode8_8C_inst0_O,Decode8_8B_inst0_O,Decode8_8A_inst0_O,Decode8_89_inst0_O,Decode8_88_inst0_O,Decode8_87_inst0_O,Decode8_86_inst0_O,Decode8_85_inst0_O,Decode8_84_inst0_O,Decode8_83_inst0_O,Decode8_82_inst0_O,Decode8_81_inst0_O,Decode8_80_inst0_O,Decode8_7F_inst0_O,Decode8_7E_inst0_O,Decode8_7D_inst0_O,Decode8_7C_inst0_O,Decode8_7B_inst0_O,Decode8_7A_inst0_O,Decode8_79_inst0_O,Decode8_78_inst0_O,Decode8_77_inst0_O,Decode8_76_inst0_O,Decode8_75_inst0_O,Decode8_74_inst0_O,Decode8_73_inst0_O,Decode8_72_inst0_O,Decode8_71_inst0_O,Decode8_70_inst0_O,Decode8_6F_inst0_O,Decode8_6E_inst0_O,Decode8_6D_inst0_O,Decode8_6C_inst0_O,Decode8_6B_inst0_O,Decode8_6A_inst0_O,Decode8_69_inst0_O,Decode8_68_inst0_O,Decode8_67_inst0_O,Decode8_66_inst0_O,Decode8_65_inst0_O,Decode8_64_inst0_O,Decode8_63_inst0_O,Decode8_62_inst0_O,Decode8_61_inst0_O,Decode8_60_inst0_O,Decode8_5F_inst0_O,Decode8_5E_inst0_O,Decode8_5D_inst0_O,Decode8_5C_inst0_O,Decode8_5B_inst0_O,Decode8_5A_inst0_O,Decode8_59_inst0_O,Decode8_58_inst0_O,Decode8_57_inst0_O,Decode8_56_inst0_O,Decode8_55_inst0_O,Decode8_54_inst0_O,Decode8_53_inst0_O,Decode8_52_inst0_O,Decode8_51_inst0_O,Decode8_50_inst0_O,Decode8_4F_inst0_O,Decode8_4E_inst0_O,Decode8_4D_inst0_O,Decode8_4C_inst0_O,Decode8_4B_inst0_O,Decode8_4A_inst0_O,Decode8_49_inst0_O,Decode8_48_inst0_O,Decode8_47_inst0_O,Decode8_46_inst0_O,Decode8_45_inst0_O,Decode8_44_inst0_O,Decode8_43_inst0_O,Decode8_42_inst0_O,Decode8_41_inst0_O,Decode8_40_inst0_O,Decode8_3F_inst0_O,Decode8_3E_inst0_O,Decode8_3D_inst0_O,Decode8_3C_inst0_O,Decode8_3B_inst0_O,Decode8_3A_inst0_O,Decode8_39_inst0_O,Decode8_38_inst0_O,Decode8_37_inst0_O,Decode8_36_inst0_O,Decode8_35_inst0_O,Decode8_34_inst0_O,Decode8_33_inst0_O,Decode8_32_inst0_O,Decode8_31_inst0_O,Decode8_30_inst0_O,Decode8_2F_inst0_O,Decode8_2E_inst0_O,Decode8_2D_inst0_O,Decode8_2C_inst0_O,Decode8_2B_inst0_O,Decode8_2A_inst0_O,Decode8_29_inst0_O,Decode8_28_inst0_O,Decode8_27_inst0_O,Decode8_26_inst0_O,Decode8_25_inst0_O,Decode8_24_inst0_O,Decode8_23_inst0_O,Decode8_22_inst0_O,Decode8_21_inst0_O,Decode8_20_inst0_O,Decode8_1F_inst0_O,Decode8_1E_inst0_O,Decode8_1D_inst0_O,Decode8_1C_inst0_O,Decode8_1B_inst0_O,Decode8_1A_inst0_O,Decode8_19_inst0_O,Decode8_18_inst0_O,Decode8_17_inst0_O,Decode8_16_inst0_O,Decode8_15_inst0_O,Decode8_14_inst0_O,Decode8_13_inst0_O,Decode8_12_inst0_O,Decode8_11_inst0_O,Decode8_10_inst0_O,Decode8_F_inst0_O,Decode8_E_inst0_O,Decode8_D_inst0_O,Decode8_C_inst0_O,Decode8_B_inst0_O,Decode8_A_inst0_O,Decode8_9_inst0_O,Decode8_8_inst0_O,Decode8_7_inst0_O,Decode8_6_inst0_O,Decode8_5_inst0_O,Decode8_4_inst0_O,Decode8_3_inst0_O,Decode8_2_inst0_O,Decode8_1_inst0_O,Decode8_0_inst0_O};
endmodule

