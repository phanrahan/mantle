module coreir_add #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 + in1;
endmodule

module coreir_add2_wrapped (
    input [1:0] I0,
    input [1:0] I1,
    output [1:0] O
);
wire [1:0] coreir_add2_inst0_in0;
wire [1:0] coreir_add2_inst0_in1;
wire [1:0] coreir_add2_inst0_out;
assign coreir_add2_inst0_in0 = I0;
assign coreir_add2_inst0_in1 = I1;
coreir_add #(
    .width(2)
) coreir_add2_inst0 (
    .in0(coreir_add2_inst0_in0),
    .in1(coreir_add2_inst0_in1),
    .out(coreir_add2_inst0_out)
);
assign O = coreir_add2_inst0_out;
endmodule

