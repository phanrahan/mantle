module FixedASR4_3 (input [3:0] I, output [3:0] O);
assign O = {I[3],I[3],I[3],I[3]};
endmodule

