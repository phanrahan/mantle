module Decode8 (input [7:0] I, output  O);
wire  LUT4_inst0_O;
wire  LUT4_inst1_O;
wire  MUXF5_inst0_O;
wire  LUT4_inst2_O;
wire  LUT4_inst3_O;
wire  MUXF5_inst1_O;
wire  MUXF6_inst0_O;
wire  LUT4_inst4_O;
wire  LUT4_inst5_O;
wire  MUXF5_inst2_O;
wire  LUT4_inst6_O;
wire  LUT4_inst7_O;
wire  MUXF5_inst3_O;
wire  MUXF6_inst1_O;
wire  MUXF7_inst0_O;
wire  LUT4_inst8_O;
wire  LUT4_inst9_O;
wire  MUXF5_inst4_O;
wire  LUT4_inst10_O;
wire  LUT4_inst11_O;
wire  MUXF5_inst5_O;
wire  MUXF6_inst2_O;
wire  LUT4_inst12_O;
wire  LUT4_inst13_O;
wire  MUXF5_inst6_O;
wire  LUT4_inst14_O;
wire  LUT4_inst15_O;
wire  MUXF5_inst7_O;
wire  MUXF6_inst3_O;
wire  MUXF7_inst1_O;
wire  MUXF8_inst0_O;
LUT4 #(.INIT(16'h0001)) LUT4_inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst1_O));
MUXF5 MUXF5_inst0 (.I0(LUT4_inst0_O), .I1(LUT4_inst1_O), .S(I[4]), .O(MUXF5_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst3_O));
MUXF5 MUXF5_inst1 (.I0(LUT4_inst2_O), .I1(LUT4_inst3_O), .S(I[4]), .O(MUXF5_inst1_O));
MUXF6 MUXF6_inst0 (.I0(MUXF5_inst0_O), .I1(MUXF5_inst1_O), .S(I[5]), .O(MUXF6_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst5_O));
MUXF5 MUXF5_inst2 (.I0(LUT4_inst4_O), .I1(LUT4_inst5_O), .S(I[4]), .O(MUXF5_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst7_O));
MUXF5 MUXF5_inst3 (.I0(LUT4_inst6_O), .I1(LUT4_inst7_O), .S(I[4]), .O(MUXF5_inst3_O));
MUXF6 MUXF6_inst1 (.I0(MUXF5_inst2_O), .I1(MUXF5_inst3_O), .S(I[5]), .O(MUXF6_inst1_O));
MUXF7 MUXF7_inst0 (.I0(MUXF6_inst0_O), .I1(MUXF6_inst1_O), .S(I[6]), .O(MUXF7_inst0_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst8_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst9_O));
MUXF5 MUXF5_inst4 (.I0(LUT4_inst8_O), .I1(LUT4_inst9_O), .S(I[4]), .O(MUXF5_inst4_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst10_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst11_O));
MUXF5 MUXF5_inst5 (.I0(LUT4_inst10_O), .I1(LUT4_inst11_O), .S(I[4]), .O(MUXF5_inst5_O));
MUXF6 MUXF6_inst2 (.I0(MUXF5_inst4_O), .I1(MUXF5_inst5_O), .S(I[5]), .O(MUXF6_inst2_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst12_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst13_O));
MUXF5 MUXF5_inst6 (.I0(LUT4_inst12_O), .I1(LUT4_inst13_O), .S(I[4]), .O(MUXF5_inst6_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst14_O));
LUT4 #(.INIT(16'h0000)) LUT4_inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(LUT4_inst15_O));
MUXF5 MUXF5_inst7 (.I0(LUT4_inst14_O), .I1(LUT4_inst15_O), .S(I[4]), .O(MUXF5_inst7_O));
MUXF6 MUXF6_inst3 (.I0(MUXF5_inst6_O), .I1(MUXF5_inst7_O), .S(I[5]), .O(MUXF6_inst3_O));
MUXF7 MUXF7_inst1 (.I0(MUXF6_inst2_O), .I1(MUXF6_inst3_O), .S(I[6]), .O(MUXF7_inst1_O));
MUXF8 MUXF8_inst0 (.I0(MUXF7_inst0_O), .I1(MUXF7_inst1_O), .S(I[7]), .O(MUXF8_inst0_O));
assign O = MUXF8_inst0_O;
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire  Decode8_inst0_O;
wire  Decode8_inst1_O;
wire  Decode8_inst2_O;
wire  Decode8_inst3_O;
wire  Decode8_inst4_O;
wire  Decode8_inst5_O;
wire  Decode8_inst6_O;
wire  Decode8_inst7_O;
wire  Decode8_inst8_O;
wire  Decode8_inst9_O;
wire  Decode8_inst10_O;
wire  Decode8_inst11_O;
wire  Decode8_inst12_O;
wire  Decode8_inst13_O;
wire  Decode8_inst14_O;
wire  Decode8_inst15_O;
wire  Decode8_inst16_O;
wire  Decode8_inst17_O;
wire  Decode8_inst18_O;
wire  Decode8_inst19_O;
wire  Decode8_inst20_O;
wire  Decode8_inst21_O;
wire  Decode8_inst22_O;
wire  Decode8_inst23_O;
wire  Decode8_inst24_O;
wire  Decode8_inst25_O;
wire  Decode8_inst26_O;
wire  Decode8_inst27_O;
wire  Decode8_inst28_O;
wire  Decode8_inst29_O;
wire  Decode8_inst30_O;
wire  Decode8_inst31_O;
wire  Decode8_inst32_O;
wire  Decode8_inst33_O;
wire  Decode8_inst34_O;
wire  Decode8_inst35_O;
wire  Decode8_inst36_O;
wire  Decode8_inst37_O;
wire  Decode8_inst38_O;
wire  Decode8_inst39_O;
wire  Decode8_inst40_O;
wire  Decode8_inst41_O;
wire  Decode8_inst42_O;
wire  Decode8_inst43_O;
wire  Decode8_inst44_O;
wire  Decode8_inst45_O;
wire  Decode8_inst46_O;
wire  Decode8_inst47_O;
wire  Decode8_inst48_O;
wire  Decode8_inst49_O;
wire  Decode8_inst50_O;
wire  Decode8_inst51_O;
wire  Decode8_inst52_O;
wire  Decode8_inst53_O;
wire  Decode8_inst54_O;
wire  Decode8_inst55_O;
wire  Decode8_inst56_O;
wire  Decode8_inst57_O;
wire  Decode8_inst58_O;
wire  Decode8_inst59_O;
wire  Decode8_inst60_O;
wire  Decode8_inst61_O;
wire  Decode8_inst62_O;
wire  Decode8_inst63_O;
wire  Decode8_inst64_O;
wire  Decode8_inst65_O;
wire  Decode8_inst66_O;
wire  Decode8_inst67_O;
wire  Decode8_inst68_O;
wire  Decode8_inst69_O;
wire  Decode8_inst70_O;
wire  Decode8_inst71_O;
wire  Decode8_inst72_O;
wire  Decode8_inst73_O;
wire  Decode8_inst74_O;
wire  Decode8_inst75_O;
wire  Decode8_inst76_O;
wire  Decode8_inst77_O;
wire  Decode8_inst78_O;
wire  Decode8_inst79_O;
wire  Decode8_inst80_O;
wire  Decode8_inst81_O;
wire  Decode8_inst82_O;
wire  Decode8_inst83_O;
wire  Decode8_inst84_O;
wire  Decode8_inst85_O;
wire  Decode8_inst86_O;
wire  Decode8_inst87_O;
wire  Decode8_inst88_O;
wire  Decode8_inst89_O;
wire  Decode8_inst90_O;
wire  Decode8_inst91_O;
wire  Decode8_inst92_O;
wire  Decode8_inst93_O;
wire  Decode8_inst94_O;
wire  Decode8_inst95_O;
wire  Decode8_inst96_O;
wire  Decode8_inst97_O;
wire  Decode8_inst98_O;
wire  Decode8_inst99_O;
wire  Decode8_inst100_O;
wire  Decode8_inst101_O;
wire  Decode8_inst102_O;
wire  Decode8_inst103_O;
wire  Decode8_inst104_O;
wire  Decode8_inst105_O;
wire  Decode8_inst106_O;
wire  Decode8_inst107_O;
wire  Decode8_inst108_O;
wire  Decode8_inst109_O;
wire  Decode8_inst110_O;
wire  Decode8_inst111_O;
wire  Decode8_inst112_O;
wire  Decode8_inst113_O;
wire  Decode8_inst114_O;
wire  Decode8_inst115_O;
wire  Decode8_inst116_O;
wire  Decode8_inst117_O;
wire  Decode8_inst118_O;
wire  Decode8_inst119_O;
wire  Decode8_inst120_O;
wire  Decode8_inst121_O;
wire  Decode8_inst122_O;
wire  Decode8_inst123_O;
wire  Decode8_inst124_O;
wire  Decode8_inst125_O;
wire  Decode8_inst126_O;
wire  Decode8_inst127_O;
wire  Decode8_inst128_O;
wire  Decode8_inst129_O;
wire  Decode8_inst130_O;
wire  Decode8_inst131_O;
wire  Decode8_inst132_O;
wire  Decode8_inst133_O;
wire  Decode8_inst134_O;
wire  Decode8_inst135_O;
wire  Decode8_inst136_O;
wire  Decode8_inst137_O;
wire  Decode8_inst138_O;
wire  Decode8_inst139_O;
wire  Decode8_inst140_O;
wire  Decode8_inst141_O;
wire  Decode8_inst142_O;
wire  Decode8_inst143_O;
wire  Decode8_inst144_O;
wire  Decode8_inst145_O;
wire  Decode8_inst146_O;
wire  Decode8_inst147_O;
wire  Decode8_inst148_O;
wire  Decode8_inst149_O;
wire  Decode8_inst150_O;
wire  Decode8_inst151_O;
wire  Decode8_inst152_O;
wire  Decode8_inst153_O;
wire  Decode8_inst154_O;
wire  Decode8_inst155_O;
wire  Decode8_inst156_O;
wire  Decode8_inst157_O;
wire  Decode8_inst158_O;
wire  Decode8_inst159_O;
wire  Decode8_inst160_O;
wire  Decode8_inst161_O;
wire  Decode8_inst162_O;
wire  Decode8_inst163_O;
wire  Decode8_inst164_O;
wire  Decode8_inst165_O;
wire  Decode8_inst166_O;
wire  Decode8_inst167_O;
wire  Decode8_inst168_O;
wire  Decode8_inst169_O;
wire  Decode8_inst170_O;
wire  Decode8_inst171_O;
wire  Decode8_inst172_O;
wire  Decode8_inst173_O;
wire  Decode8_inst174_O;
wire  Decode8_inst175_O;
wire  Decode8_inst176_O;
wire  Decode8_inst177_O;
wire  Decode8_inst178_O;
wire  Decode8_inst179_O;
wire  Decode8_inst180_O;
wire  Decode8_inst181_O;
wire  Decode8_inst182_O;
wire  Decode8_inst183_O;
wire  Decode8_inst184_O;
wire  Decode8_inst185_O;
wire  Decode8_inst186_O;
wire  Decode8_inst187_O;
wire  Decode8_inst188_O;
wire  Decode8_inst189_O;
wire  Decode8_inst190_O;
wire  Decode8_inst191_O;
wire  Decode8_inst192_O;
wire  Decode8_inst193_O;
wire  Decode8_inst194_O;
wire  Decode8_inst195_O;
wire  Decode8_inst196_O;
wire  Decode8_inst197_O;
wire  Decode8_inst198_O;
wire  Decode8_inst199_O;
wire  Decode8_inst200_O;
wire  Decode8_inst201_O;
wire  Decode8_inst202_O;
wire  Decode8_inst203_O;
wire  Decode8_inst204_O;
wire  Decode8_inst205_O;
wire  Decode8_inst206_O;
wire  Decode8_inst207_O;
wire  Decode8_inst208_O;
wire  Decode8_inst209_O;
wire  Decode8_inst210_O;
wire  Decode8_inst211_O;
wire  Decode8_inst212_O;
wire  Decode8_inst213_O;
wire  Decode8_inst214_O;
wire  Decode8_inst215_O;
wire  Decode8_inst216_O;
wire  Decode8_inst217_O;
wire  Decode8_inst218_O;
wire  Decode8_inst219_O;
wire  Decode8_inst220_O;
wire  Decode8_inst221_O;
wire  Decode8_inst222_O;
wire  Decode8_inst223_O;
wire  Decode8_inst224_O;
wire  Decode8_inst225_O;
wire  Decode8_inst226_O;
wire  Decode8_inst227_O;
wire  Decode8_inst228_O;
wire  Decode8_inst229_O;
wire  Decode8_inst230_O;
wire  Decode8_inst231_O;
wire  Decode8_inst232_O;
wire  Decode8_inst233_O;
wire  Decode8_inst234_O;
wire  Decode8_inst235_O;
wire  Decode8_inst236_O;
wire  Decode8_inst237_O;
wire  Decode8_inst238_O;
wire  Decode8_inst239_O;
wire  Decode8_inst240_O;
wire  Decode8_inst241_O;
wire  Decode8_inst242_O;
wire  Decode8_inst243_O;
wire  Decode8_inst244_O;
wire  Decode8_inst245_O;
wire  Decode8_inst246_O;
wire  Decode8_inst247_O;
wire  Decode8_inst248_O;
wire  Decode8_inst249_O;
wire  Decode8_inst250_O;
wire  Decode8_inst251_O;
wire  Decode8_inst252_O;
wire  Decode8_inst253_O;
wire  Decode8_inst254_O;
wire  Decode8_inst255_O;
Decode8 Decode8_inst0 (.I(I), .O(Decode8_inst0_O));
Decode8 Decode8_inst1 (.I(I), .O(Decode8_inst1_O));
Decode8 Decode8_inst2 (.I(I), .O(Decode8_inst2_O));
Decode8 Decode8_inst3 (.I(I), .O(Decode8_inst3_O));
Decode8 Decode8_inst4 (.I(I), .O(Decode8_inst4_O));
Decode8 Decode8_inst5 (.I(I), .O(Decode8_inst5_O));
Decode8 Decode8_inst6 (.I(I), .O(Decode8_inst6_O));
Decode8 Decode8_inst7 (.I(I), .O(Decode8_inst7_O));
Decode8 Decode8_inst8 (.I(I), .O(Decode8_inst8_O));
Decode8 Decode8_inst9 (.I(I), .O(Decode8_inst9_O));
Decode8 Decode8_inst10 (.I(I), .O(Decode8_inst10_O));
Decode8 Decode8_inst11 (.I(I), .O(Decode8_inst11_O));
Decode8 Decode8_inst12 (.I(I), .O(Decode8_inst12_O));
Decode8 Decode8_inst13 (.I(I), .O(Decode8_inst13_O));
Decode8 Decode8_inst14 (.I(I), .O(Decode8_inst14_O));
Decode8 Decode8_inst15 (.I(I), .O(Decode8_inst15_O));
Decode8 Decode8_inst16 (.I(I), .O(Decode8_inst16_O));
Decode8 Decode8_inst17 (.I(I), .O(Decode8_inst17_O));
Decode8 Decode8_inst18 (.I(I), .O(Decode8_inst18_O));
Decode8 Decode8_inst19 (.I(I), .O(Decode8_inst19_O));
Decode8 Decode8_inst20 (.I(I), .O(Decode8_inst20_O));
Decode8 Decode8_inst21 (.I(I), .O(Decode8_inst21_O));
Decode8 Decode8_inst22 (.I(I), .O(Decode8_inst22_O));
Decode8 Decode8_inst23 (.I(I), .O(Decode8_inst23_O));
Decode8 Decode8_inst24 (.I(I), .O(Decode8_inst24_O));
Decode8 Decode8_inst25 (.I(I), .O(Decode8_inst25_O));
Decode8 Decode8_inst26 (.I(I), .O(Decode8_inst26_O));
Decode8 Decode8_inst27 (.I(I), .O(Decode8_inst27_O));
Decode8 Decode8_inst28 (.I(I), .O(Decode8_inst28_O));
Decode8 Decode8_inst29 (.I(I), .O(Decode8_inst29_O));
Decode8 Decode8_inst30 (.I(I), .O(Decode8_inst30_O));
Decode8 Decode8_inst31 (.I(I), .O(Decode8_inst31_O));
Decode8 Decode8_inst32 (.I(I), .O(Decode8_inst32_O));
Decode8 Decode8_inst33 (.I(I), .O(Decode8_inst33_O));
Decode8 Decode8_inst34 (.I(I), .O(Decode8_inst34_O));
Decode8 Decode8_inst35 (.I(I), .O(Decode8_inst35_O));
Decode8 Decode8_inst36 (.I(I), .O(Decode8_inst36_O));
Decode8 Decode8_inst37 (.I(I), .O(Decode8_inst37_O));
Decode8 Decode8_inst38 (.I(I), .O(Decode8_inst38_O));
Decode8 Decode8_inst39 (.I(I), .O(Decode8_inst39_O));
Decode8 Decode8_inst40 (.I(I), .O(Decode8_inst40_O));
Decode8 Decode8_inst41 (.I(I), .O(Decode8_inst41_O));
Decode8 Decode8_inst42 (.I(I), .O(Decode8_inst42_O));
Decode8 Decode8_inst43 (.I(I), .O(Decode8_inst43_O));
Decode8 Decode8_inst44 (.I(I), .O(Decode8_inst44_O));
Decode8 Decode8_inst45 (.I(I), .O(Decode8_inst45_O));
Decode8 Decode8_inst46 (.I(I), .O(Decode8_inst46_O));
Decode8 Decode8_inst47 (.I(I), .O(Decode8_inst47_O));
Decode8 Decode8_inst48 (.I(I), .O(Decode8_inst48_O));
Decode8 Decode8_inst49 (.I(I), .O(Decode8_inst49_O));
Decode8 Decode8_inst50 (.I(I), .O(Decode8_inst50_O));
Decode8 Decode8_inst51 (.I(I), .O(Decode8_inst51_O));
Decode8 Decode8_inst52 (.I(I), .O(Decode8_inst52_O));
Decode8 Decode8_inst53 (.I(I), .O(Decode8_inst53_O));
Decode8 Decode8_inst54 (.I(I), .O(Decode8_inst54_O));
Decode8 Decode8_inst55 (.I(I), .O(Decode8_inst55_O));
Decode8 Decode8_inst56 (.I(I), .O(Decode8_inst56_O));
Decode8 Decode8_inst57 (.I(I), .O(Decode8_inst57_O));
Decode8 Decode8_inst58 (.I(I), .O(Decode8_inst58_O));
Decode8 Decode8_inst59 (.I(I), .O(Decode8_inst59_O));
Decode8 Decode8_inst60 (.I(I), .O(Decode8_inst60_O));
Decode8 Decode8_inst61 (.I(I), .O(Decode8_inst61_O));
Decode8 Decode8_inst62 (.I(I), .O(Decode8_inst62_O));
Decode8 Decode8_inst63 (.I(I), .O(Decode8_inst63_O));
Decode8 Decode8_inst64 (.I(I), .O(Decode8_inst64_O));
Decode8 Decode8_inst65 (.I(I), .O(Decode8_inst65_O));
Decode8 Decode8_inst66 (.I(I), .O(Decode8_inst66_O));
Decode8 Decode8_inst67 (.I(I), .O(Decode8_inst67_O));
Decode8 Decode8_inst68 (.I(I), .O(Decode8_inst68_O));
Decode8 Decode8_inst69 (.I(I), .O(Decode8_inst69_O));
Decode8 Decode8_inst70 (.I(I), .O(Decode8_inst70_O));
Decode8 Decode8_inst71 (.I(I), .O(Decode8_inst71_O));
Decode8 Decode8_inst72 (.I(I), .O(Decode8_inst72_O));
Decode8 Decode8_inst73 (.I(I), .O(Decode8_inst73_O));
Decode8 Decode8_inst74 (.I(I), .O(Decode8_inst74_O));
Decode8 Decode8_inst75 (.I(I), .O(Decode8_inst75_O));
Decode8 Decode8_inst76 (.I(I), .O(Decode8_inst76_O));
Decode8 Decode8_inst77 (.I(I), .O(Decode8_inst77_O));
Decode8 Decode8_inst78 (.I(I), .O(Decode8_inst78_O));
Decode8 Decode8_inst79 (.I(I), .O(Decode8_inst79_O));
Decode8 Decode8_inst80 (.I(I), .O(Decode8_inst80_O));
Decode8 Decode8_inst81 (.I(I), .O(Decode8_inst81_O));
Decode8 Decode8_inst82 (.I(I), .O(Decode8_inst82_O));
Decode8 Decode8_inst83 (.I(I), .O(Decode8_inst83_O));
Decode8 Decode8_inst84 (.I(I), .O(Decode8_inst84_O));
Decode8 Decode8_inst85 (.I(I), .O(Decode8_inst85_O));
Decode8 Decode8_inst86 (.I(I), .O(Decode8_inst86_O));
Decode8 Decode8_inst87 (.I(I), .O(Decode8_inst87_O));
Decode8 Decode8_inst88 (.I(I), .O(Decode8_inst88_O));
Decode8 Decode8_inst89 (.I(I), .O(Decode8_inst89_O));
Decode8 Decode8_inst90 (.I(I), .O(Decode8_inst90_O));
Decode8 Decode8_inst91 (.I(I), .O(Decode8_inst91_O));
Decode8 Decode8_inst92 (.I(I), .O(Decode8_inst92_O));
Decode8 Decode8_inst93 (.I(I), .O(Decode8_inst93_O));
Decode8 Decode8_inst94 (.I(I), .O(Decode8_inst94_O));
Decode8 Decode8_inst95 (.I(I), .O(Decode8_inst95_O));
Decode8 Decode8_inst96 (.I(I), .O(Decode8_inst96_O));
Decode8 Decode8_inst97 (.I(I), .O(Decode8_inst97_O));
Decode8 Decode8_inst98 (.I(I), .O(Decode8_inst98_O));
Decode8 Decode8_inst99 (.I(I), .O(Decode8_inst99_O));
Decode8 Decode8_inst100 (.I(I), .O(Decode8_inst100_O));
Decode8 Decode8_inst101 (.I(I), .O(Decode8_inst101_O));
Decode8 Decode8_inst102 (.I(I), .O(Decode8_inst102_O));
Decode8 Decode8_inst103 (.I(I), .O(Decode8_inst103_O));
Decode8 Decode8_inst104 (.I(I), .O(Decode8_inst104_O));
Decode8 Decode8_inst105 (.I(I), .O(Decode8_inst105_O));
Decode8 Decode8_inst106 (.I(I), .O(Decode8_inst106_O));
Decode8 Decode8_inst107 (.I(I), .O(Decode8_inst107_O));
Decode8 Decode8_inst108 (.I(I), .O(Decode8_inst108_O));
Decode8 Decode8_inst109 (.I(I), .O(Decode8_inst109_O));
Decode8 Decode8_inst110 (.I(I), .O(Decode8_inst110_O));
Decode8 Decode8_inst111 (.I(I), .O(Decode8_inst111_O));
Decode8 Decode8_inst112 (.I(I), .O(Decode8_inst112_O));
Decode8 Decode8_inst113 (.I(I), .O(Decode8_inst113_O));
Decode8 Decode8_inst114 (.I(I), .O(Decode8_inst114_O));
Decode8 Decode8_inst115 (.I(I), .O(Decode8_inst115_O));
Decode8 Decode8_inst116 (.I(I), .O(Decode8_inst116_O));
Decode8 Decode8_inst117 (.I(I), .O(Decode8_inst117_O));
Decode8 Decode8_inst118 (.I(I), .O(Decode8_inst118_O));
Decode8 Decode8_inst119 (.I(I), .O(Decode8_inst119_O));
Decode8 Decode8_inst120 (.I(I), .O(Decode8_inst120_O));
Decode8 Decode8_inst121 (.I(I), .O(Decode8_inst121_O));
Decode8 Decode8_inst122 (.I(I), .O(Decode8_inst122_O));
Decode8 Decode8_inst123 (.I(I), .O(Decode8_inst123_O));
Decode8 Decode8_inst124 (.I(I), .O(Decode8_inst124_O));
Decode8 Decode8_inst125 (.I(I), .O(Decode8_inst125_O));
Decode8 Decode8_inst126 (.I(I), .O(Decode8_inst126_O));
Decode8 Decode8_inst127 (.I(I), .O(Decode8_inst127_O));
Decode8 Decode8_inst128 (.I(I), .O(Decode8_inst128_O));
Decode8 Decode8_inst129 (.I(I), .O(Decode8_inst129_O));
Decode8 Decode8_inst130 (.I(I), .O(Decode8_inst130_O));
Decode8 Decode8_inst131 (.I(I), .O(Decode8_inst131_O));
Decode8 Decode8_inst132 (.I(I), .O(Decode8_inst132_O));
Decode8 Decode8_inst133 (.I(I), .O(Decode8_inst133_O));
Decode8 Decode8_inst134 (.I(I), .O(Decode8_inst134_O));
Decode8 Decode8_inst135 (.I(I), .O(Decode8_inst135_O));
Decode8 Decode8_inst136 (.I(I), .O(Decode8_inst136_O));
Decode8 Decode8_inst137 (.I(I), .O(Decode8_inst137_O));
Decode8 Decode8_inst138 (.I(I), .O(Decode8_inst138_O));
Decode8 Decode8_inst139 (.I(I), .O(Decode8_inst139_O));
Decode8 Decode8_inst140 (.I(I), .O(Decode8_inst140_O));
Decode8 Decode8_inst141 (.I(I), .O(Decode8_inst141_O));
Decode8 Decode8_inst142 (.I(I), .O(Decode8_inst142_O));
Decode8 Decode8_inst143 (.I(I), .O(Decode8_inst143_O));
Decode8 Decode8_inst144 (.I(I), .O(Decode8_inst144_O));
Decode8 Decode8_inst145 (.I(I), .O(Decode8_inst145_O));
Decode8 Decode8_inst146 (.I(I), .O(Decode8_inst146_O));
Decode8 Decode8_inst147 (.I(I), .O(Decode8_inst147_O));
Decode8 Decode8_inst148 (.I(I), .O(Decode8_inst148_O));
Decode8 Decode8_inst149 (.I(I), .O(Decode8_inst149_O));
Decode8 Decode8_inst150 (.I(I), .O(Decode8_inst150_O));
Decode8 Decode8_inst151 (.I(I), .O(Decode8_inst151_O));
Decode8 Decode8_inst152 (.I(I), .O(Decode8_inst152_O));
Decode8 Decode8_inst153 (.I(I), .O(Decode8_inst153_O));
Decode8 Decode8_inst154 (.I(I), .O(Decode8_inst154_O));
Decode8 Decode8_inst155 (.I(I), .O(Decode8_inst155_O));
Decode8 Decode8_inst156 (.I(I), .O(Decode8_inst156_O));
Decode8 Decode8_inst157 (.I(I), .O(Decode8_inst157_O));
Decode8 Decode8_inst158 (.I(I), .O(Decode8_inst158_O));
Decode8 Decode8_inst159 (.I(I), .O(Decode8_inst159_O));
Decode8 Decode8_inst160 (.I(I), .O(Decode8_inst160_O));
Decode8 Decode8_inst161 (.I(I), .O(Decode8_inst161_O));
Decode8 Decode8_inst162 (.I(I), .O(Decode8_inst162_O));
Decode8 Decode8_inst163 (.I(I), .O(Decode8_inst163_O));
Decode8 Decode8_inst164 (.I(I), .O(Decode8_inst164_O));
Decode8 Decode8_inst165 (.I(I), .O(Decode8_inst165_O));
Decode8 Decode8_inst166 (.I(I), .O(Decode8_inst166_O));
Decode8 Decode8_inst167 (.I(I), .O(Decode8_inst167_O));
Decode8 Decode8_inst168 (.I(I), .O(Decode8_inst168_O));
Decode8 Decode8_inst169 (.I(I), .O(Decode8_inst169_O));
Decode8 Decode8_inst170 (.I(I), .O(Decode8_inst170_O));
Decode8 Decode8_inst171 (.I(I), .O(Decode8_inst171_O));
Decode8 Decode8_inst172 (.I(I), .O(Decode8_inst172_O));
Decode8 Decode8_inst173 (.I(I), .O(Decode8_inst173_O));
Decode8 Decode8_inst174 (.I(I), .O(Decode8_inst174_O));
Decode8 Decode8_inst175 (.I(I), .O(Decode8_inst175_O));
Decode8 Decode8_inst176 (.I(I), .O(Decode8_inst176_O));
Decode8 Decode8_inst177 (.I(I), .O(Decode8_inst177_O));
Decode8 Decode8_inst178 (.I(I), .O(Decode8_inst178_O));
Decode8 Decode8_inst179 (.I(I), .O(Decode8_inst179_O));
Decode8 Decode8_inst180 (.I(I), .O(Decode8_inst180_O));
Decode8 Decode8_inst181 (.I(I), .O(Decode8_inst181_O));
Decode8 Decode8_inst182 (.I(I), .O(Decode8_inst182_O));
Decode8 Decode8_inst183 (.I(I), .O(Decode8_inst183_O));
Decode8 Decode8_inst184 (.I(I), .O(Decode8_inst184_O));
Decode8 Decode8_inst185 (.I(I), .O(Decode8_inst185_O));
Decode8 Decode8_inst186 (.I(I), .O(Decode8_inst186_O));
Decode8 Decode8_inst187 (.I(I), .O(Decode8_inst187_O));
Decode8 Decode8_inst188 (.I(I), .O(Decode8_inst188_O));
Decode8 Decode8_inst189 (.I(I), .O(Decode8_inst189_O));
Decode8 Decode8_inst190 (.I(I), .O(Decode8_inst190_O));
Decode8 Decode8_inst191 (.I(I), .O(Decode8_inst191_O));
Decode8 Decode8_inst192 (.I(I), .O(Decode8_inst192_O));
Decode8 Decode8_inst193 (.I(I), .O(Decode8_inst193_O));
Decode8 Decode8_inst194 (.I(I), .O(Decode8_inst194_O));
Decode8 Decode8_inst195 (.I(I), .O(Decode8_inst195_O));
Decode8 Decode8_inst196 (.I(I), .O(Decode8_inst196_O));
Decode8 Decode8_inst197 (.I(I), .O(Decode8_inst197_O));
Decode8 Decode8_inst198 (.I(I), .O(Decode8_inst198_O));
Decode8 Decode8_inst199 (.I(I), .O(Decode8_inst199_O));
Decode8 Decode8_inst200 (.I(I), .O(Decode8_inst200_O));
Decode8 Decode8_inst201 (.I(I), .O(Decode8_inst201_O));
Decode8 Decode8_inst202 (.I(I), .O(Decode8_inst202_O));
Decode8 Decode8_inst203 (.I(I), .O(Decode8_inst203_O));
Decode8 Decode8_inst204 (.I(I), .O(Decode8_inst204_O));
Decode8 Decode8_inst205 (.I(I), .O(Decode8_inst205_O));
Decode8 Decode8_inst206 (.I(I), .O(Decode8_inst206_O));
Decode8 Decode8_inst207 (.I(I), .O(Decode8_inst207_O));
Decode8 Decode8_inst208 (.I(I), .O(Decode8_inst208_O));
Decode8 Decode8_inst209 (.I(I), .O(Decode8_inst209_O));
Decode8 Decode8_inst210 (.I(I), .O(Decode8_inst210_O));
Decode8 Decode8_inst211 (.I(I), .O(Decode8_inst211_O));
Decode8 Decode8_inst212 (.I(I), .O(Decode8_inst212_O));
Decode8 Decode8_inst213 (.I(I), .O(Decode8_inst213_O));
Decode8 Decode8_inst214 (.I(I), .O(Decode8_inst214_O));
Decode8 Decode8_inst215 (.I(I), .O(Decode8_inst215_O));
Decode8 Decode8_inst216 (.I(I), .O(Decode8_inst216_O));
Decode8 Decode8_inst217 (.I(I), .O(Decode8_inst217_O));
Decode8 Decode8_inst218 (.I(I), .O(Decode8_inst218_O));
Decode8 Decode8_inst219 (.I(I), .O(Decode8_inst219_O));
Decode8 Decode8_inst220 (.I(I), .O(Decode8_inst220_O));
Decode8 Decode8_inst221 (.I(I), .O(Decode8_inst221_O));
Decode8 Decode8_inst222 (.I(I), .O(Decode8_inst222_O));
Decode8 Decode8_inst223 (.I(I), .O(Decode8_inst223_O));
Decode8 Decode8_inst224 (.I(I), .O(Decode8_inst224_O));
Decode8 Decode8_inst225 (.I(I), .O(Decode8_inst225_O));
Decode8 Decode8_inst226 (.I(I), .O(Decode8_inst226_O));
Decode8 Decode8_inst227 (.I(I), .O(Decode8_inst227_O));
Decode8 Decode8_inst228 (.I(I), .O(Decode8_inst228_O));
Decode8 Decode8_inst229 (.I(I), .O(Decode8_inst229_O));
Decode8 Decode8_inst230 (.I(I), .O(Decode8_inst230_O));
Decode8 Decode8_inst231 (.I(I), .O(Decode8_inst231_O));
Decode8 Decode8_inst232 (.I(I), .O(Decode8_inst232_O));
Decode8 Decode8_inst233 (.I(I), .O(Decode8_inst233_O));
Decode8 Decode8_inst234 (.I(I), .O(Decode8_inst234_O));
Decode8 Decode8_inst235 (.I(I), .O(Decode8_inst235_O));
Decode8 Decode8_inst236 (.I(I), .O(Decode8_inst236_O));
Decode8 Decode8_inst237 (.I(I), .O(Decode8_inst237_O));
Decode8 Decode8_inst238 (.I(I), .O(Decode8_inst238_O));
Decode8 Decode8_inst239 (.I(I), .O(Decode8_inst239_O));
Decode8 Decode8_inst240 (.I(I), .O(Decode8_inst240_O));
Decode8 Decode8_inst241 (.I(I), .O(Decode8_inst241_O));
Decode8 Decode8_inst242 (.I(I), .O(Decode8_inst242_O));
Decode8 Decode8_inst243 (.I(I), .O(Decode8_inst243_O));
Decode8 Decode8_inst244 (.I(I), .O(Decode8_inst244_O));
Decode8 Decode8_inst245 (.I(I), .O(Decode8_inst245_O));
Decode8 Decode8_inst246 (.I(I), .O(Decode8_inst246_O));
Decode8 Decode8_inst247 (.I(I), .O(Decode8_inst247_O));
Decode8 Decode8_inst248 (.I(I), .O(Decode8_inst248_O));
Decode8 Decode8_inst249 (.I(I), .O(Decode8_inst249_O));
Decode8 Decode8_inst250 (.I(I), .O(Decode8_inst250_O));
Decode8 Decode8_inst251 (.I(I), .O(Decode8_inst251_O));
Decode8 Decode8_inst252 (.I(I), .O(Decode8_inst252_O));
Decode8 Decode8_inst253 (.I(I), .O(Decode8_inst253_O));
Decode8 Decode8_inst254 (.I(I), .O(Decode8_inst254_O));
Decode8 Decode8_inst255 (.I(I), .O(Decode8_inst255_O));
assign O = {Decode8_inst255_O,Decode8_inst254_O,Decode8_inst253_O,Decode8_inst252_O,Decode8_inst251_O,Decode8_inst250_O,Decode8_inst249_O,Decode8_inst248_O,Decode8_inst247_O,Decode8_inst246_O,Decode8_inst245_O,Decode8_inst244_O,Decode8_inst243_O,Decode8_inst242_O,Decode8_inst241_O,Decode8_inst240_O,Decode8_inst239_O,Decode8_inst238_O,Decode8_inst237_O,Decode8_inst236_O,Decode8_inst235_O,Decode8_inst234_O,Decode8_inst233_O,Decode8_inst232_O,Decode8_inst231_O,Decode8_inst230_O,Decode8_inst229_O,Decode8_inst228_O,Decode8_inst227_O,Decode8_inst226_O,Decode8_inst225_O,Decode8_inst224_O,Decode8_inst223_O,Decode8_inst222_O,Decode8_inst221_O,Decode8_inst220_O,Decode8_inst219_O,Decode8_inst218_O,Decode8_inst217_O,Decode8_inst216_O,Decode8_inst215_O,Decode8_inst214_O,Decode8_inst213_O,Decode8_inst212_O,Decode8_inst211_O,Decode8_inst210_O,Decode8_inst209_O,Decode8_inst208_O,Decode8_inst207_O,Decode8_inst206_O,Decode8_inst205_O,Decode8_inst204_O,Decode8_inst203_O,Decode8_inst202_O,Decode8_inst201_O,Decode8_inst200_O,Decode8_inst199_O,Decode8_inst198_O,Decode8_inst197_O,Decode8_inst196_O,Decode8_inst195_O,Decode8_inst194_O,Decode8_inst193_O,Decode8_inst192_O,Decode8_inst191_O,Decode8_inst190_O,Decode8_inst189_O,Decode8_inst188_O,Decode8_inst187_O,Decode8_inst186_O,Decode8_inst185_O,Decode8_inst184_O,Decode8_inst183_O,Decode8_inst182_O,Decode8_inst181_O,Decode8_inst180_O,Decode8_inst179_O,Decode8_inst178_O,Decode8_inst177_O,Decode8_inst176_O,Decode8_inst175_O,Decode8_inst174_O,Decode8_inst173_O,Decode8_inst172_O,Decode8_inst171_O,Decode8_inst170_O,Decode8_inst169_O,Decode8_inst168_O,Decode8_inst167_O,Decode8_inst166_O,Decode8_inst165_O,Decode8_inst164_O,Decode8_inst163_O,Decode8_inst162_O,Decode8_inst161_O,Decode8_inst160_O,Decode8_inst159_O,Decode8_inst158_O,Decode8_inst157_O,Decode8_inst156_O,Decode8_inst155_O,Decode8_inst154_O,Decode8_inst153_O,Decode8_inst152_O,Decode8_inst151_O,Decode8_inst150_O,Decode8_inst149_O,Decode8_inst148_O,Decode8_inst147_O,Decode8_inst146_O,Decode8_inst145_O,Decode8_inst144_O,Decode8_inst143_O,Decode8_inst142_O,Decode8_inst141_O,Decode8_inst140_O,Decode8_inst139_O,Decode8_inst138_O,Decode8_inst137_O,Decode8_inst136_O,Decode8_inst135_O,Decode8_inst134_O,Decode8_inst133_O,Decode8_inst132_O,Decode8_inst131_O,Decode8_inst130_O,Decode8_inst129_O,Decode8_inst128_O,Decode8_inst127_O,Decode8_inst126_O,Decode8_inst125_O,Decode8_inst124_O,Decode8_inst123_O,Decode8_inst122_O,Decode8_inst121_O,Decode8_inst120_O,Decode8_inst119_O,Decode8_inst118_O,Decode8_inst117_O,Decode8_inst116_O,Decode8_inst115_O,Decode8_inst114_O,Decode8_inst113_O,Decode8_inst112_O,Decode8_inst111_O,Decode8_inst110_O,Decode8_inst109_O,Decode8_inst108_O,Decode8_inst107_O,Decode8_inst106_O,Decode8_inst105_O,Decode8_inst104_O,Decode8_inst103_O,Decode8_inst102_O,Decode8_inst101_O,Decode8_inst100_O,Decode8_inst99_O,Decode8_inst98_O,Decode8_inst97_O,Decode8_inst96_O,Decode8_inst95_O,Decode8_inst94_O,Decode8_inst93_O,Decode8_inst92_O,Decode8_inst91_O,Decode8_inst90_O,Decode8_inst89_O,Decode8_inst88_O,Decode8_inst87_O,Decode8_inst86_O,Decode8_inst85_O,Decode8_inst84_O,Decode8_inst83_O,Decode8_inst82_O,Decode8_inst81_O,Decode8_inst80_O,Decode8_inst79_O,Decode8_inst78_O,Decode8_inst77_O,Decode8_inst76_O,Decode8_inst75_O,Decode8_inst74_O,Decode8_inst73_O,Decode8_inst72_O,Decode8_inst71_O,Decode8_inst70_O,Decode8_inst69_O,Decode8_inst68_O,Decode8_inst67_O,Decode8_inst66_O,Decode8_inst65_O,Decode8_inst64_O,Decode8_inst63_O,Decode8_inst62_O,Decode8_inst61_O,Decode8_inst60_O,Decode8_inst59_O,Decode8_inst58_O,Decode8_inst57_O,Decode8_inst56_O,Decode8_inst55_O,Decode8_inst54_O,Decode8_inst53_O,Decode8_inst52_O,Decode8_inst51_O,Decode8_inst50_O,Decode8_inst49_O,Decode8_inst48_O,Decode8_inst47_O,Decode8_inst46_O,Decode8_inst45_O,Decode8_inst44_O,Decode8_inst43_O,Decode8_inst42_O,Decode8_inst41_O,Decode8_inst40_O,Decode8_inst39_O,Decode8_inst38_O,Decode8_inst37_O,Decode8_inst36_O,Decode8_inst35_O,Decode8_inst34_O,Decode8_inst33_O,Decode8_inst32_O,Decode8_inst31_O,Decode8_inst30_O,Decode8_inst29_O,Decode8_inst28_O,Decode8_inst27_O,Decode8_inst26_O,Decode8_inst25_O,Decode8_inst24_O,Decode8_inst23_O,Decode8_inst22_O,Decode8_inst21_O,Decode8_inst20_O,Decode8_inst19_O,Decode8_inst18_O,Decode8_inst17_O,Decode8_inst16_O,Decode8_inst15_O,Decode8_inst14_O,Decode8_inst13_O,Decode8_inst12_O,Decode8_inst11_O,Decode8_inst10_O,Decode8_inst9_O,Decode8_inst8_O,Decode8_inst7_O,Decode8_inst6_O,Decode8_inst5_O,Decode8_inst4_O,Decode8_inst3_O,Decode8_inst2_O,Decode8_inst1_O,Decode8_inst0_O};
endmodule

