module main (output [7:0] LED, input  CLKIN, input [7:0] SWITCH);
wire [15:0] inst0_DO;
wire [1:0] inst0_DOP;
RAMB16_S18 #(.INIT_39(256'h9F009E009D009C009B009A009900980097009600950094009300920091009000),
.INIT_2A(256'hAF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A000),
.INIT_2B(256'hBF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B000),
.INIT_2C(256'hCF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C000),
.INIT_2D(256'hDF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D000),
.INIT_2E(256'hEF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E000),
.INIT_2F(256'hFF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F000),
.INIT_0B(256'hBF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B000),
.INIT_0C(256'hCF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C000),
.INIT_0A(256'hAF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A000),
.INIT_0F(256'hFF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F000),
.INIT_0D(256'hDF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D000),
.INIT_0E(256'hEF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E000),
.WRITE_MODE("WRITE_FIRST"),
.INIT_15(256'h5F005E005D005C005B005A005900580057005600550054005300520051005000),
.INIT_14(256'h4F004E004D004C004B004A004900480047004600450044004300420041004000),
.INIT_17(256'h7F007E007D007C007B007A007900780077007600750074007300720071007000),
.INIT_16(256'h6F006E006D006C006B006A006900680067006600650064006300620061006000),
.INIT_11(256'h1F001E001D001C001B001A001900180017001600150014001300120011001000),
.INIT_10(256'h0F000E000D000C000B000A000900080007000600050004000300020001000000),
.INIT_13(256'h3F003E003D003C003B003A003900380037003600350034003300320031003000),
.INIT_12(256'h2F002E002D002C002B002A002900280027002600250024002300220021002000),
.INIT_19(256'h9F009E009D009C009B009A009900980097009600950094009300920091009000),
.INIT_18(256'h8F008E008D008C008B008A008900880087008600850084008300820081008000),
.INIT(16'h0000),
.INIT_38(256'h8F008E008D008C008B008A008900880087008600850084008300820081008000),
.INIT_33(256'h3F003E003D003C003B003A003900380037003600350034003300320031003000),
.INIT_32(256'h2F002E002D002C002B002A002900280027002600250024002300220021002000),
.INIT_31(256'h1F001E001D001C001B001A001900180017001600150014001300120011001000),
.INIT_30(256'h0F000E000D000C000B000A000900080007000600050004000300020001000000),
.INIT_37(256'h7F007E007D007C007B007A007900780077007600750074007300720071007000),
.INIT_36(256'h6F006E006D006C006B006A006900680067006600650064006300620061006000),
.INIT_35(256'h5F005E005D005C005B005A005900580057005600550054005300520051005000),
.INIT_34(256'h4F004E004D004C004B004A004900480047004600450044004300420041004000),
.SRVAL(16'h0000),
.INIT_3C(256'hCF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C000),
.INIT_3B(256'hBF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B000),
.INIT_3A(256'hAF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A000),
.INIT_3F(256'hFF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F000),
.INIT_3E(256'hEF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E000),
.INIT_3D(256'hDF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D000),
.INIT_1E(256'hEF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E000),
.INIT_1D(256'hDF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D000),
.INIT_1F(256'hFF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F000),
.INIT_1A(256'hAF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A000),
.INIT_1C(256'hCF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C000),
.INIT_1B(256'hBF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B000),
.INIT_02(256'h2F002E002D002C002B002A002900280027002600250024002300220021002000),
.INIT_03(256'h3F003E003D003C003B003A003900380037003600350034003300320031003000),
.INIT_00(256'h0F000E000D000C000B000A000900080007000600050004000300020001000000),
.INIT_01(256'h1F001E001D001C001B001A001900180017001600150014001300120011001000),
.INIT_06(256'h6F006E006D006C006B006A006900680067006600650064006300620061006000),
.INIT_07(256'h7F007E007D007C007B007A007900780077007600750074007300720071007000),
.INIT_04(256'h4F004E004D004C004B004A004900480047004600450044004300420041004000),
.INIT_05(256'h5F005E005D005C005B005A005900580057005600550054005300520051005000),
.INIT_08(256'h8F008E008D008C008B008A008900880087008600850084008300820081008000),
.INIT_09(256'h9F009E009D009C009B009A009900980097009600950094009300920091009000),
.INIT_28(256'h8F008E008D008C008B008A008900880087008600850084008300820081008000),
.INIT_29(256'h9F009E009D009C009B009A009900980097009600950094009300920091009000),
.INIT_20(256'h0F000E000D000C000B000A000900080007000600050004000300020001000000),
.INIT_21(256'h1F001E001D001C001B001A001900180017001600150014001300120011001000),
.INIT_22(256'h2F002E002D002C002B002A002900280027002600250024002300220021002000),
.INIT_23(256'h3F003E003D003C003B003A003900380037003600350034003300320031003000),
.INIT_24(256'h4F004E004D004C004B004A004900480047004600450044004300420041004000),
.INIT_25(256'h5F005E005D005C005B005A005900580057005600550054005300520051005000),
.INIT_26(256'h6F006E006D006C006B006A006900680067006600650064006300620061006000),
.INIT_27(256'h7F007E007D007C007B007A007900780077007600750074007300720071007000)) inst0 (.DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .DIP({1'b0,1'b0}), .DO(inst0_DO), .DOP(inst0_DOP), .ADDR({1'b0,1'b0,SWITCH[7],SWITCH[6],SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .CLK(CLKIN), .EN(1'b1), .SSR(1'b0), .WE(1'b0));
assign LED = {inst0_DO[15],inst0_DO[14],inst0_DO[13],inst0_DO[12],inst0_DO[11],inst0_DO[10],inst0_DO[9],inst0_DO[8]};
endmodule

