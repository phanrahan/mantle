module main (output [7:0] LED, input  CLKIN, input [7:0] SWITCH);
wire [15:0] inst0_DO;
wire [1:0] inst0_DOP;
RAMB16_S18 #(.INIT_39(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_2A(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_2B(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_2C(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_2D(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_2E(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_2F(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_0B(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_0C(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_0A(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_0F(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_0D(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_0E(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.WRITE_MODE("WRITE_FIRST"),
.INIT_15(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_14(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_17(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_16(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_11(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_10(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_13(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_12(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_19(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_18(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT(18'h00000),
.INIT_38(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
.INIT_32(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
.INITP_02(256'h5555555555555555555555555555555500000000000000000000000000000000),
.INIT_37(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_36(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_35(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_34(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_05(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.SRVAL(18'h00000),
.INIT_3C(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_3B(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_3A(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_01(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_3F(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_3E(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_3D(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_1E(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_33(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_1F(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_1A(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INITP_00(256'h5555555555555555555555555555555500000000000000000000000000000000),
.INIT_1C(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_1B(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_31(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_02(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_03(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_00(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_30(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_06(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_07(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_04(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_1D(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INITP_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
.INIT_08(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_09(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INITP_04(256'h5555555555555555555555555555555500000000000000000000000000000000),
.INIT_28(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_29(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INITP_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
.INIT_23(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000),
.INIT_20(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_21(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_22(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INITP_06(256'h5555555555555555555555555555555500000000000000000000000000000000),
.INIT_24(256'h3C003800340030002C002800240020001C001800140010000C00080004000000),
.INIT_25(256'h7C007800740070006C006800640060005C005800540050004C00480044004000),
.INIT_26(256'hBC00B800B400B000AC00A800A400A0009C009800940090008C00880084008000),
.INIT_27(256'hFC00F800F400F000EC00E800E400E000DC00D800D400D000CC00C800C400C000)) inst0 (.DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .DIP({1'b0,1'b0}), .DO(inst0_DO), .DOP(inst0_DOP), .ADDR({1'b0,1'b0,SWITCH[7],SWITCH[6],SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .CLK(CLKIN), .EN(1'b1), .SSR(1'b0), .WE(1'b0));
assign LED = {inst0_DOP[1],inst0_DOP[0],inst0_DO[15],inst0_DO[14],inst0_DO[13],inst0_DO[12],inst0_DO[11],inst0_DO[10]};
endmodule

