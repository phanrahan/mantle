module coreir_eq #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output out);
  assign out = in0 == in1;
endmodule

module Decode998 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h63), .out(O));
endmodule

module Decode988 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h62), .out(O));
endmodule

module Decode98 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h09), .out(O));
endmodule

module Decode978 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h61), .out(O));
endmodule

module Decode968 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h60), .out(O));
endmodule

module Decode958 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5f), .out(O));
endmodule

module Decode948 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5e), .out(O));
endmodule

module Decode938 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5d), .out(O));
endmodule

module Decode928 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5c), .out(O));
endmodule

module Decode918 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5b), .out(O));
endmodule

module Decode908 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h5a), .out(O));
endmodule

module Decode898 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h59), .out(O));
endmodule

module Decode888 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h58), .out(O));
endmodule

module Decode88 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h08), .out(O));
endmodule

module Decode878 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h57), .out(O));
endmodule

module Decode868 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h56), .out(O));
endmodule

module Decode858 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h55), .out(O));
endmodule

module Decode848 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h54), .out(O));
endmodule

module Decode838 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h53), .out(O));
endmodule

module Decode828 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h52), .out(O));
endmodule

module Decode818 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h51), .out(O));
endmodule

module Decode808 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h50), .out(O));
endmodule

module Decode798 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4f), .out(O));
endmodule

module Decode788 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4e), .out(O));
endmodule

module Decode78 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h07), .out(O));
endmodule

module Decode778 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4d), .out(O));
endmodule

module Decode768 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4c), .out(O));
endmodule

module Decode758 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4b), .out(O));
endmodule

module Decode748 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h4a), .out(O));
endmodule

module Decode738 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h49), .out(O));
endmodule

module Decode728 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h48), .out(O));
endmodule

module Decode718 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h47), .out(O));
endmodule

module Decode708 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h46), .out(O));
endmodule

module Decode698 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h45), .out(O));
endmodule

module Decode688 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h44), .out(O));
endmodule

module Decode68 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h06), .out(O));
endmodule

module Decode678 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h43), .out(O));
endmodule

module Decode668 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h42), .out(O));
endmodule

module Decode658 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h41), .out(O));
endmodule

module Decode648 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h40), .out(O));
endmodule

module Decode638 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3f), .out(O));
endmodule

module Decode628 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3e), .out(O));
endmodule

module Decode618 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3d), .out(O));
endmodule

module Decode608 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3c), .out(O));
endmodule

module Decode598 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3b), .out(O));
endmodule

module Decode588 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h3a), .out(O));
endmodule

module Decode58 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h05), .out(O));
endmodule

module Decode578 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h39), .out(O));
endmodule

module Decode568 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h38), .out(O));
endmodule

module Decode558 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h37), .out(O));
endmodule

module Decode548 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h36), .out(O));
endmodule

module Decode538 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h35), .out(O));
endmodule

module Decode528 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h34), .out(O));
endmodule

module Decode518 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h33), .out(O));
endmodule

module Decode508 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h32), .out(O));
endmodule

module Decode498 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h31), .out(O));
endmodule

module Decode488 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h30), .out(O));
endmodule

module Decode48 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h04), .out(O));
endmodule

module Decode478 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2f), .out(O));
endmodule

module Decode468 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2e), .out(O));
endmodule

module Decode458 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2d), .out(O));
endmodule

module Decode448 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2c), .out(O));
endmodule

module Decode438 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2b), .out(O));
endmodule

module Decode428 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h2a), .out(O));
endmodule

module Decode418 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h29), .out(O));
endmodule

module Decode408 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h28), .out(O));
endmodule

module Decode398 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h27), .out(O));
endmodule

module Decode388 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h26), .out(O));
endmodule

module Decode38 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h03), .out(O));
endmodule

module Decode378 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h25), .out(O));
endmodule

module Decode368 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h24), .out(O));
endmodule

module Decode358 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h23), .out(O));
endmodule

module Decode348 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h22), .out(O));
endmodule

module Decode338 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h21), .out(O));
endmodule

module Decode328 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h20), .out(O));
endmodule

module Decode318 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1f), .out(O));
endmodule

module Decode308 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1e), .out(O));
endmodule

module Decode298 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1d), .out(O));
endmodule

module Decode288 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1c), .out(O));
endmodule

module Decode28 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h02), .out(O));
endmodule

module Decode278 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1b), .out(O));
endmodule

module Decode268 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h1a), .out(O));
endmodule

module Decode258 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h19), .out(O));
endmodule

module Decode2558 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hff), .out(O));
endmodule

module Decode2548 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hfe), .out(O));
endmodule

module Decode2538 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hfd), .out(O));
endmodule

module Decode2528 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hfc), .out(O));
endmodule

module Decode2518 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hfb), .out(O));
endmodule

module Decode2508 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hfa), .out(O));
endmodule

module Decode2498 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf9), .out(O));
endmodule

module Decode2488 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf8), .out(O));
endmodule

module Decode248 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h18), .out(O));
endmodule

module Decode2478 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf7), .out(O));
endmodule

module Decode2468 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf6), .out(O));
endmodule

module Decode2458 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf5), .out(O));
endmodule

module Decode2448 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf4), .out(O));
endmodule

module Decode2438 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf3), .out(O));
endmodule

module Decode2428 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf2), .out(O));
endmodule

module Decode2418 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf1), .out(O));
endmodule

module Decode2408 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hf0), .out(O));
endmodule

module Decode2398 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hef), .out(O));
endmodule

module Decode2388 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hee), .out(O));
endmodule

module Decode238 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h17), .out(O));
endmodule

module Decode2378 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hed), .out(O));
endmodule

module Decode2368 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hec), .out(O));
endmodule

module Decode2358 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'heb), .out(O));
endmodule

module Decode2348 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hea), .out(O));
endmodule

module Decode2338 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he9), .out(O));
endmodule

module Decode2328 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he8), .out(O));
endmodule

module Decode2318 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he7), .out(O));
endmodule

module Decode2308 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he6), .out(O));
endmodule

module Decode2298 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he5), .out(O));
endmodule

module Decode2288 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he4), .out(O));
endmodule

module Decode228 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h16), .out(O));
endmodule

module Decode2278 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he3), .out(O));
endmodule

module Decode2268 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he2), .out(O));
endmodule

module Decode2258 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he1), .out(O));
endmodule

module Decode2248 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'he0), .out(O));
endmodule

module Decode2238 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hdf), .out(O));
endmodule

module Decode2228 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hde), .out(O));
endmodule

module Decode2218 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hdd), .out(O));
endmodule

module Decode2208 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hdc), .out(O));
endmodule

module Decode2198 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hdb), .out(O));
endmodule

module Decode2188 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hda), .out(O));
endmodule

module Decode218 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h15), .out(O));
endmodule

module Decode2178 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd9), .out(O));
endmodule

module Decode2168 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd8), .out(O));
endmodule

module Decode2158 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd7), .out(O));
endmodule

module Decode2148 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd6), .out(O));
endmodule

module Decode2138 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd5), .out(O));
endmodule

module Decode2128 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd4), .out(O));
endmodule

module Decode2118 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd3), .out(O));
endmodule

module Decode2108 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd2), .out(O));
endmodule

module Decode2098 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd1), .out(O));
endmodule

module Decode2088 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hd0), .out(O));
endmodule

module Decode208 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h14), .out(O));
endmodule

module Decode2078 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hcf), .out(O));
endmodule

module Decode2068 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hce), .out(O));
endmodule

module Decode2058 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hcd), .out(O));
endmodule

module Decode2048 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hcc), .out(O));
endmodule

module Decode2038 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hcb), .out(O));
endmodule

module Decode2028 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hca), .out(O));
endmodule

module Decode2018 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc9), .out(O));
endmodule

module Decode2008 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc8), .out(O));
endmodule

module Decode1998 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc7), .out(O));
endmodule

module Decode1988 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc6), .out(O));
endmodule

module Decode198 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h13), .out(O));
endmodule

module Decode1978 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc5), .out(O));
endmodule

module Decode1968 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc4), .out(O));
endmodule

module Decode1958 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc3), .out(O));
endmodule

module Decode1948 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc2), .out(O));
endmodule

module Decode1938 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc1), .out(O));
endmodule

module Decode1928 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hc0), .out(O));
endmodule

module Decode1918 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hbf), .out(O));
endmodule

module Decode1908 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hbe), .out(O));
endmodule

module Decode1898 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hbd), .out(O));
endmodule

module Decode1888 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hbc), .out(O));
endmodule

module Decode188 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h12), .out(O));
endmodule

module Decode1878 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hbb), .out(O));
endmodule

module Decode1868 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hba), .out(O));
endmodule

module Decode1858 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb9), .out(O));
endmodule

module Decode1848 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb8), .out(O));
endmodule

module Decode1838 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb7), .out(O));
endmodule

module Decode1828 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb6), .out(O));
endmodule

module Decode1818 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb5), .out(O));
endmodule

module Decode1808 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb4), .out(O));
endmodule

module Decode18 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h01), .out(O));
endmodule

module Decode1798 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb3), .out(O));
endmodule

module Decode1788 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb2), .out(O));
endmodule

module Decode178 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h11), .out(O));
endmodule

module Decode1778 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb1), .out(O));
endmodule

module Decode1768 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hb0), .out(O));
endmodule

module Decode1758 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'haf), .out(O));
endmodule

module Decode1748 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hae), .out(O));
endmodule

module Decode1738 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'had), .out(O));
endmodule

module Decode1728 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hac), .out(O));
endmodule

module Decode1718 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'hab), .out(O));
endmodule

module Decode1708 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'haa), .out(O));
endmodule

module Decode1698 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha9), .out(O));
endmodule

module Decode1688 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha8), .out(O));
endmodule

module Decode168 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h10), .out(O));
endmodule

module Decode1678 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha7), .out(O));
endmodule

module Decode1668 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha6), .out(O));
endmodule

module Decode1658 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha5), .out(O));
endmodule

module Decode1648 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha4), .out(O));
endmodule

module Decode1638 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha3), .out(O));
endmodule

module Decode1628 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha2), .out(O));
endmodule

module Decode1618 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha1), .out(O));
endmodule

module Decode1608 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'ha0), .out(O));
endmodule

module Decode1598 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9f), .out(O));
endmodule

module Decode1588 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9e), .out(O));
endmodule

module Decode158 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0f), .out(O));
endmodule

module Decode1578 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9d), .out(O));
endmodule

module Decode1568 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9c), .out(O));
endmodule

module Decode1558 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9b), .out(O));
endmodule

module Decode1548 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h9a), .out(O));
endmodule

module Decode1538 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h99), .out(O));
endmodule

module Decode1528 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h98), .out(O));
endmodule

module Decode1518 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h97), .out(O));
endmodule

module Decode1508 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h96), .out(O));
endmodule

module Decode1498 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h95), .out(O));
endmodule

module Decode1488 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h94), .out(O));
endmodule

module Decode148 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0e), .out(O));
endmodule

module Decode1478 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h93), .out(O));
endmodule

module Decode1468 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h92), .out(O));
endmodule

module Decode1458 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h91), .out(O));
endmodule

module Decode1448 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h90), .out(O));
endmodule

module Decode1438 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8f), .out(O));
endmodule

module Decode1428 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8e), .out(O));
endmodule

module Decode1418 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8d), .out(O));
endmodule

module Decode1408 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8c), .out(O));
endmodule

module Decode1398 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8b), .out(O));
endmodule

module Decode1388 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h8a), .out(O));
endmodule

module Decode138 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0d), .out(O));
endmodule

module Decode1378 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h89), .out(O));
endmodule

module Decode1368 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h88), .out(O));
endmodule

module Decode1358 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h87), .out(O));
endmodule

module Decode1348 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h86), .out(O));
endmodule

module Decode1338 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h85), .out(O));
endmodule

module Decode1328 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h84), .out(O));
endmodule

module Decode1318 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h83), .out(O));
endmodule

module Decode1308 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h82), .out(O));
endmodule

module Decode1298 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h81), .out(O));
endmodule

module Decode1288 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h80), .out(O));
endmodule

module Decode128 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0c), .out(O));
endmodule

module Decode1278 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7f), .out(O));
endmodule

module Decode1268 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7e), .out(O));
endmodule

module Decode1258 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7d), .out(O));
endmodule

module Decode1248 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7c), .out(O));
endmodule

module Decode1238 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7b), .out(O));
endmodule

module Decode1228 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h7a), .out(O));
endmodule

module Decode1218 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h79), .out(O));
endmodule

module Decode1208 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h78), .out(O));
endmodule

module Decode1198 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h77), .out(O));
endmodule

module Decode1188 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h76), .out(O));
endmodule

module Decode118 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0b), .out(O));
endmodule

module Decode1178 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h75), .out(O));
endmodule

module Decode1168 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h74), .out(O));
endmodule

module Decode1158 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h73), .out(O));
endmodule

module Decode1148 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h72), .out(O));
endmodule

module Decode1138 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h71), .out(O));
endmodule

module Decode1128 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h70), .out(O));
endmodule

module Decode1118 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6f), .out(O));
endmodule

module Decode1108 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6e), .out(O));
endmodule

module Decode1098 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6d), .out(O));
endmodule

module Decode1088 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6c), .out(O));
endmodule

module Decode108 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h0a), .out(O));
endmodule

module Decode1078 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6b), .out(O));
endmodule

module Decode1068 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h6a), .out(O));
endmodule

module Decode1058 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h69), .out(O));
endmodule

module Decode1048 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h68), .out(O));
endmodule

module Decode1038 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h67), .out(O));
endmodule

module Decode1028 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h66), .out(O));
endmodule

module Decode1018 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h65), .out(O));
endmodule

module Decode1008 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h64), .out(O));
endmodule

module Decode08 (input [7:0] I, output O);
coreir_eq #(.width(8)) coreir_eq_8_inst0(.in0(I), .in1(8'h00), .out(O));
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire Decode08_inst0_O;
wire Decode1008_inst0_O;
wire Decode1018_inst0_O;
wire Decode1028_inst0_O;
wire Decode1038_inst0_O;
wire Decode1048_inst0_O;
wire Decode1058_inst0_O;
wire Decode1068_inst0_O;
wire Decode1078_inst0_O;
wire Decode1088_inst0_O;
wire Decode108_inst0_O;
wire Decode1098_inst0_O;
wire Decode1108_inst0_O;
wire Decode1118_inst0_O;
wire Decode1128_inst0_O;
wire Decode1138_inst0_O;
wire Decode1148_inst0_O;
wire Decode1158_inst0_O;
wire Decode1168_inst0_O;
wire Decode1178_inst0_O;
wire Decode1188_inst0_O;
wire Decode118_inst0_O;
wire Decode1198_inst0_O;
wire Decode1208_inst0_O;
wire Decode1218_inst0_O;
wire Decode1228_inst0_O;
wire Decode1238_inst0_O;
wire Decode1248_inst0_O;
wire Decode1258_inst0_O;
wire Decode1268_inst0_O;
wire Decode1278_inst0_O;
wire Decode1288_inst0_O;
wire Decode128_inst0_O;
wire Decode1298_inst0_O;
wire Decode1308_inst0_O;
wire Decode1318_inst0_O;
wire Decode1328_inst0_O;
wire Decode1338_inst0_O;
wire Decode1348_inst0_O;
wire Decode1358_inst0_O;
wire Decode1368_inst0_O;
wire Decode1378_inst0_O;
wire Decode1388_inst0_O;
wire Decode138_inst0_O;
wire Decode1398_inst0_O;
wire Decode1408_inst0_O;
wire Decode1418_inst0_O;
wire Decode1428_inst0_O;
wire Decode1438_inst0_O;
wire Decode1448_inst0_O;
wire Decode1458_inst0_O;
wire Decode1468_inst0_O;
wire Decode1478_inst0_O;
wire Decode1488_inst0_O;
wire Decode148_inst0_O;
wire Decode1498_inst0_O;
wire Decode1508_inst0_O;
wire Decode1518_inst0_O;
wire Decode1528_inst0_O;
wire Decode1538_inst0_O;
wire Decode1548_inst0_O;
wire Decode1558_inst0_O;
wire Decode1568_inst0_O;
wire Decode1578_inst0_O;
wire Decode1588_inst0_O;
wire Decode158_inst0_O;
wire Decode1598_inst0_O;
wire Decode1608_inst0_O;
wire Decode1618_inst0_O;
wire Decode1628_inst0_O;
wire Decode1638_inst0_O;
wire Decode1648_inst0_O;
wire Decode1658_inst0_O;
wire Decode1668_inst0_O;
wire Decode1678_inst0_O;
wire Decode1688_inst0_O;
wire Decode168_inst0_O;
wire Decode1698_inst0_O;
wire Decode1708_inst0_O;
wire Decode1718_inst0_O;
wire Decode1728_inst0_O;
wire Decode1738_inst0_O;
wire Decode1748_inst0_O;
wire Decode1758_inst0_O;
wire Decode1768_inst0_O;
wire Decode1778_inst0_O;
wire Decode1788_inst0_O;
wire Decode178_inst0_O;
wire Decode1798_inst0_O;
wire Decode1808_inst0_O;
wire Decode1818_inst0_O;
wire Decode1828_inst0_O;
wire Decode1838_inst0_O;
wire Decode1848_inst0_O;
wire Decode1858_inst0_O;
wire Decode1868_inst0_O;
wire Decode1878_inst0_O;
wire Decode1888_inst0_O;
wire Decode188_inst0_O;
wire Decode1898_inst0_O;
wire Decode18_inst0_O;
wire Decode1908_inst0_O;
wire Decode1918_inst0_O;
wire Decode1928_inst0_O;
wire Decode1938_inst0_O;
wire Decode1948_inst0_O;
wire Decode1958_inst0_O;
wire Decode1968_inst0_O;
wire Decode1978_inst0_O;
wire Decode1988_inst0_O;
wire Decode198_inst0_O;
wire Decode1998_inst0_O;
wire Decode2008_inst0_O;
wire Decode2018_inst0_O;
wire Decode2028_inst0_O;
wire Decode2038_inst0_O;
wire Decode2048_inst0_O;
wire Decode2058_inst0_O;
wire Decode2068_inst0_O;
wire Decode2078_inst0_O;
wire Decode2088_inst0_O;
wire Decode208_inst0_O;
wire Decode2098_inst0_O;
wire Decode2108_inst0_O;
wire Decode2118_inst0_O;
wire Decode2128_inst0_O;
wire Decode2138_inst0_O;
wire Decode2148_inst0_O;
wire Decode2158_inst0_O;
wire Decode2168_inst0_O;
wire Decode2178_inst0_O;
wire Decode2188_inst0_O;
wire Decode218_inst0_O;
wire Decode2198_inst0_O;
wire Decode2208_inst0_O;
wire Decode2218_inst0_O;
wire Decode2228_inst0_O;
wire Decode2238_inst0_O;
wire Decode2248_inst0_O;
wire Decode2258_inst0_O;
wire Decode2268_inst0_O;
wire Decode2278_inst0_O;
wire Decode2288_inst0_O;
wire Decode228_inst0_O;
wire Decode2298_inst0_O;
wire Decode2308_inst0_O;
wire Decode2318_inst0_O;
wire Decode2328_inst0_O;
wire Decode2338_inst0_O;
wire Decode2348_inst0_O;
wire Decode2358_inst0_O;
wire Decode2368_inst0_O;
wire Decode2378_inst0_O;
wire Decode2388_inst0_O;
wire Decode238_inst0_O;
wire Decode2398_inst0_O;
wire Decode2408_inst0_O;
wire Decode2418_inst0_O;
wire Decode2428_inst0_O;
wire Decode2438_inst0_O;
wire Decode2448_inst0_O;
wire Decode2458_inst0_O;
wire Decode2468_inst0_O;
wire Decode2478_inst0_O;
wire Decode2488_inst0_O;
wire Decode248_inst0_O;
wire Decode2498_inst0_O;
wire Decode2508_inst0_O;
wire Decode2518_inst0_O;
wire Decode2528_inst0_O;
wire Decode2538_inst0_O;
wire Decode2548_inst0_O;
wire Decode2558_inst0_O;
wire Decode258_inst0_O;
wire Decode268_inst0_O;
wire Decode278_inst0_O;
wire Decode288_inst0_O;
wire Decode28_inst0_O;
wire Decode298_inst0_O;
wire Decode308_inst0_O;
wire Decode318_inst0_O;
wire Decode328_inst0_O;
wire Decode338_inst0_O;
wire Decode348_inst0_O;
wire Decode358_inst0_O;
wire Decode368_inst0_O;
wire Decode378_inst0_O;
wire Decode388_inst0_O;
wire Decode38_inst0_O;
wire Decode398_inst0_O;
wire Decode408_inst0_O;
wire Decode418_inst0_O;
wire Decode428_inst0_O;
wire Decode438_inst0_O;
wire Decode448_inst0_O;
wire Decode458_inst0_O;
wire Decode468_inst0_O;
wire Decode478_inst0_O;
wire Decode488_inst0_O;
wire Decode48_inst0_O;
wire Decode498_inst0_O;
wire Decode508_inst0_O;
wire Decode518_inst0_O;
wire Decode528_inst0_O;
wire Decode538_inst0_O;
wire Decode548_inst0_O;
wire Decode558_inst0_O;
wire Decode568_inst0_O;
wire Decode578_inst0_O;
wire Decode588_inst0_O;
wire Decode58_inst0_O;
wire Decode598_inst0_O;
wire Decode608_inst0_O;
wire Decode618_inst0_O;
wire Decode628_inst0_O;
wire Decode638_inst0_O;
wire Decode648_inst0_O;
wire Decode658_inst0_O;
wire Decode668_inst0_O;
wire Decode678_inst0_O;
wire Decode688_inst0_O;
wire Decode68_inst0_O;
wire Decode698_inst0_O;
wire Decode708_inst0_O;
wire Decode718_inst0_O;
wire Decode728_inst0_O;
wire Decode738_inst0_O;
wire Decode748_inst0_O;
wire Decode758_inst0_O;
wire Decode768_inst0_O;
wire Decode778_inst0_O;
wire Decode788_inst0_O;
wire Decode78_inst0_O;
wire Decode798_inst0_O;
wire Decode808_inst0_O;
wire Decode818_inst0_O;
wire Decode828_inst0_O;
wire Decode838_inst0_O;
wire Decode848_inst0_O;
wire Decode858_inst0_O;
wire Decode868_inst0_O;
wire Decode878_inst0_O;
wire Decode888_inst0_O;
wire Decode88_inst0_O;
wire Decode898_inst0_O;
wire Decode908_inst0_O;
wire Decode918_inst0_O;
wire Decode928_inst0_O;
wire Decode938_inst0_O;
wire Decode948_inst0_O;
wire Decode958_inst0_O;
wire Decode968_inst0_O;
wire Decode978_inst0_O;
wire Decode988_inst0_O;
wire Decode98_inst0_O;
wire Decode998_inst0_O;
Decode08 Decode08_inst0(.I(I), .O(Decode08_inst0_O));
Decode1008 Decode1008_inst0(.I(I), .O(Decode1008_inst0_O));
Decode1018 Decode1018_inst0(.I(I), .O(Decode1018_inst0_O));
Decode1028 Decode1028_inst0(.I(I), .O(Decode1028_inst0_O));
Decode1038 Decode1038_inst0(.I(I), .O(Decode1038_inst0_O));
Decode1048 Decode1048_inst0(.I(I), .O(Decode1048_inst0_O));
Decode1058 Decode1058_inst0(.I(I), .O(Decode1058_inst0_O));
Decode1068 Decode1068_inst0(.I(I), .O(Decode1068_inst0_O));
Decode1078 Decode1078_inst0(.I(I), .O(Decode1078_inst0_O));
Decode1088 Decode1088_inst0(.I(I), .O(Decode1088_inst0_O));
Decode108 Decode108_inst0(.I(I), .O(Decode108_inst0_O));
Decode1098 Decode1098_inst0(.I(I), .O(Decode1098_inst0_O));
Decode1108 Decode1108_inst0(.I(I), .O(Decode1108_inst0_O));
Decode1118 Decode1118_inst0(.I(I), .O(Decode1118_inst0_O));
Decode1128 Decode1128_inst0(.I(I), .O(Decode1128_inst0_O));
Decode1138 Decode1138_inst0(.I(I), .O(Decode1138_inst0_O));
Decode1148 Decode1148_inst0(.I(I), .O(Decode1148_inst0_O));
Decode1158 Decode1158_inst0(.I(I), .O(Decode1158_inst0_O));
Decode1168 Decode1168_inst0(.I(I), .O(Decode1168_inst0_O));
Decode1178 Decode1178_inst0(.I(I), .O(Decode1178_inst0_O));
Decode1188 Decode1188_inst0(.I(I), .O(Decode1188_inst0_O));
Decode118 Decode118_inst0(.I(I), .O(Decode118_inst0_O));
Decode1198 Decode1198_inst0(.I(I), .O(Decode1198_inst0_O));
Decode1208 Decode1208_inst0(.I(I), .O(Decode1208_inst0_O));
Decode1218 Decode1218_inst0(.I(I), .O(Decode1218_inst0_O));
Decode1228 Decode1228_inst0(.I(I), .O(Decode1228_inst0_O));
Decode1238 Decode1238_inst0(.I(I), .O(Decode1238_inst0_O));
Decode1248 Decode1248_inst0(.I(I), .O(Decode1248_inst0_O));
Decode1258 Decode1258_inst0(.I(I), .O(Decode1258_inst0_O));
Decode1268 Decode1268_inst0(.I(I), .O(Decode1268_inst0_O));
Decode1278 Decode1278_inst0(.I(I), .O(Decode1278_inst0_O));
Decode1288 Decode1288_inst0(.I(I), .O(Decode1288_inst0_O));
Decode128 Decode128_inst0(.I(I), .O(Decode128_inst0_O));
Decode1298 Decode1298_inst0(.I(I), .O(Decode1298_inst0_O));
Decode1308 Decode1308_inst0(.I(I), .O(Decode1308_inst0_O));
Decode1318 Decode1318_inst0(.I(I), .O(Decode1318_inst0_O));
Decode1328 Decode1328_inst0(.I(I), .O(Decode1328_inst0_O));
Decode1338 Decode1338_inst0(.I(I), .O(Decode1338_inst0_O));
Decode1348 Decode1348_inst0(.I(I), .O(Decode1348_inst0_O));
Decode1358 Decode1358_inst0(.I(I), .O(Decode1358_inst0_O));
Decode1368 Decode1368_inst0(.I(I), .O(Decode1368_inst0_O));
Decode1378 Decode1378_inst0(.I(I), .O(Decode1378_inst0_O));
Decode1388 Decode1388_inst0(.I(I), .O(Decode1388_inst0_O));
Decode138 Decode138_inst0(.I(I), .O(Decode138_inst0_O));
Decode1398 Decode1398_inst0(.I(I), .O(Decode1398_inst0_O));
Decode1408 Decode1408_inst0(.I(I), .O(Decode1408_inst0_O));
Decode1418 Decode1418_inst0(.I(I), .O(Decode1418_inst0_O));
Decode1428 Decode1428_inst0(.I(I), .O(Decode1428_inst0_O));
Decode1438 Decode1438_inst0(.I(I), .O(Decode1438_inst0_O));
Decode1448 Decode1448_inst0(.I(I), .O(Decode1448_inst0_O));
Decode1458 Decode1458_inst0(.I(I), .O(Decode1458_inst0_O));
Decode1468 Decode1468_inst0(.I(I), .O(Decode1468_inst0_O));
Decode1478 Decode1478_inst0(.I(I), .O(Decode1478_inst0_O));
Decode1488 Decode1488_inst0(.I(I), .O(Decode1488_inst0_O));
Decode148 Decode148_inst0(.I(I), .O(Decode148_inst0_O));
Decode1498 Decode1498_inst0(.I(I), .O(Decode1498_inst0_O));
Decode1508 Decode1508_inst0(.I(I), .O(Decode1508_inst0_O));
Decode1518 Decode1518_inst0(.I(I), .O(Decode1518_inst0_O));
Decode1528 Decode1528_inst0(.I(I), .O(Decode1528_inst0_O));
Decode1538 Decode1538_inst0(.I(I), .O(Decode1538_inst0_O));
Decode1548 Decode1548_inst0(.I(I), .O(Decode1548_inst0_O));
Decode1558 Decode1558_inst0(.I(I), .O(Decode1558_inst0_O));
Decode1568 Decode1568_inst0(.I(I), .O(Decode1568_inst0_O));
Decode1578 Decode1578_inst0(.I(I), .O(Decode1578_inst0_O));
Decode1588 Decode1588_inst0(.I(I), .O(Decode1588_inst0_O));
Decode158 Decode158_inst0(.I(I), .O(Decode158_inst0_O));
Decode1598 Decode1598_inst0(.I(I), .O(Decode1598_inst0_O));
Decode1608 Decode1608_inst0(.I(I), .O(Decode1608_inst0_O));
Decode1618 Decode1618_inst0(.I(I), .O(Decode1618_inst0_O));
Decode1628 Decode1628_inst0(.I(I), .O(Decode1628_inst0_O));
Decode1638 Decode1638_inst0(.I(I), .O(Decode1638_inst0_O));
Decode1648 Decode1648_inst0(.I(I), .O(Decode1648_inst0_O));
Decode1658 Decode1658_inst0(.I(I), .O(Decode1658_inst0_O));
Decode1668 Decode1668_inst0(.I(I), .O(Decode1668_inst0_O));
Decode1678 Decode1678_inst0(.I(I), .O(Decode1678_inst0_O));
Decode1688 Decode1688_inst0(.I(I), .O(Decode1688_inst0_O));
Decode168 Decode168_inst0(.I(I), .O(Decode168_inst0_O));
Decode1698 Decode1698_inst0(.I(I), .O(Decode1698_inst0_O));
Decode1708 Decode1708_inst0(.I(I), .O(Decode1708_inst0_O));
Decode1718 Decode1718_inst0(.I(I), .O(Decode1718_inst0_O));
Decode1728 Decode1728_inst0(.I(I), .O(Decode1728_inst0_O));
Decode1738 Decode1738_inst0(.I(I), .O(Decode1738_inst0_O));
Decode1748 Decode1748_inst0(.I(I), .O(Decode1748_inst0_O));
Decode1758 Decode1758_inst0(.I(I), .O(Decode1758_inst0_O));
Decode1768 Decode1768_inst0(.I(I), .O(Decode1768_inst0_O));
Decode1778 Decode1778_inst0(.I(I), .O(Decode1778_inst0_O));
Decode1788 Decode1788_inst0(.I(I), .O(Decode1788_inst0_O));
Decode178 Decode178_inst0(.I(I), .O(Decode178_inst0_O));
Decode1798 Decode1798_inst0(.I(I), .O(Decode1798_inst0_O));
Decode1808 Decode1808_inst0(.I(I), .O(Decode1808_inst0_O));
Decode1818 Decode1818_inst0(.I(I), .O(Decode1818_inst0_O));
Decode1828 Decode1828_inst0(.I(I), .O(Decode1828_inst0_O));
Decode1838 Decode1838_inst0(.I(I), .O(Decode1838_inst0_O));
Decode1848 Decode1848_inst0(.I(I), .O(Decode1848_inst0_O));
Decode1858 Decode1858_inst0(.I(I), .O(Decode1858_inst0_O));
Decode1868 Decode1868_inst0(.I(I), .O(Decode1868_inst0_O));
Decode1878 Decode1878_inst0(.I(I), .O(Decode1878_inst0_O));
Decode1888 Decode1888_inst0(.I(I), .O(Decode1888_inst0_O));
Decode188 Decode188_inst0(.I(I), .O(Decode188_inst0_O));
Decode1898 Decode1898_inst0(.I(I), .O(Decode1898_inst0_O));
Decode18 Decode18_inst0(.I(I), .O(Decode18_inst0_O));
Decode1908 Decode1908_inst0(.I(I), .O(Decode1908_inst0_O));
Decode1918 Decode1918_inst0(.I(I), .O(Decode1918_inst0_O));
Decode1928 Decode1928_inst0(.I(I), .O(Decode1928_inst0_O));
Decode1938 Decode1938_inst0(.I(I), .O(Decode1938_inst0_O));
Decode1948 Decode1948_inst0(.I(I), .O(Decode1948_inst0_O));
Decode1958 Decode1958_inst0(.I(I), .O(Decode1958_inst0_O));
Decode1968 Decode1968_inst0(.I(I), .O(Decode1968_inst0_O));
Decode1978 Decode1978_inst0(.I(I), .O(Decode1978_inst0_O));
Decode1988 Decode1988_inst0(.I(I), .O(Decode1988_inst0_O));
Decode198 Decode198_inst0(.I(I), .O(Decode198_inst0_O));
Decode1998 Decode1998_inst0(.I(I), .O(Decode1998_inst0_O));
Decode2008 Decode2008_inst0(.I(I), .O(Decode2008_inst0_O));
Decode2018 Decode2018_inst0(.I(I), .O(Decode2018_inst0_O));
Decode2028 Decode2028_inst0(.I(I), .O(Decode2028_inst0_O));
Decode2038 Decode2038_inst0(.I(I), .O(Decode2038_inst0_O));
Decode2048 Decode2048_inst0(.I(I), .O(Decode2048_inst0_O));
Decode2058 Decode2058_inst0(.I(I), .O(Decode2058_inst0_O));
Decode2068 Decode2068_inst0(.I(I), .O(Decode2068_inst0_O));
Decode2078 Decode2078_inst0(.I(I), .O(Decode2078_inst0_O));
Decode2088 Decode2088_inst0(.I(I), .O(Decode2088_inst0_O));
Decode208 Decode208_inst0(.I(I), .O(Decode208_inst0_O));
Decode2098 Decode2098_inst0(.I(I), .O(Decode2098_inst0_O));
Decode2108 Decode2108_inst0(.I(I), .O(Decode2108_inst0_O));
Decode2118 Decode2118_inst0(.I(I), .O(Decode2118_inst0_O));
Decode2128 Decode2128_inst0(.I(I), .O(Decode2128_inst0_O));
Decode2138 Decode2138_inst0(.I(I), .O(Decode2138_inst0_O));
Decode2148 Decode2148_inst0(.I(I), .O(Decode2148_inst0_O));
Decode2158 Decode2158_inst0(.I(I), .O(Decode2158_inst0_O));
Decode2168 Decode2168_inst0(.I(I), .O(Decode2168_inst0_O));
Decode2178 Decode2178_inst0(.I(I), .O(Decode2178_inst0_O));
Decode2188 Decode2188_inst0(.I(I), .O(Decode2188_inst0_O));
Decode218 Decode218_inst0(.I(I), .O(Decode218_inst0_O));
Decode2198 Decode2198_inst0(.I(I), .O(Decode2198_inst0_O));
Decode2208 Decode2208_inst0(.I(I), .O(Decode2208_inst0_O));
Decode2218 Decode2218_inst0(.I(I), .O(Decode2218_inst0_O));
Decode2228 Decode2228_inst0(.I(I), .O(Decode2228_inst0_O));
Decode2238 Decode2238_inst0(.I(I), .O(Decode2238_inst0_O));
Decode2248 Decode2248_inst0(.I(I), .O(Decode2248_inst0_O));
Decode2258 Decode2258_inst0(.I(I), .O(Decode2258_inst0_O));
Decode2268 Decode2268_inst0(.I(I), .O(Decode2268_inst0_O));
Decode2278 Decode2278_inst0(.I(I), .O(Decode2278_inst0_O));
Decode2288 Decode2288_inst0(.I(I), .O(Decode2288_inst0_O));
Decode228 Decode228_inst0(.I(I), .O(Decode228_inst0_O));
Decode2298 Decode2298_inst0(.I(I), .O(Decode2298_inst0_O));
Decode2308 Decode2308_inst0(.I(I), .O(Decode2308_inst0_O));
Decode2318 Decode2318_inst0(.I(I), .O(Decode2318_inst0_O));
Decode2328 Decode2328_inst0(.I(I), .O(Decode2328_inst0_O));
Decode2338 Decode2338_inst0(.I(I), .O(Decode2338_inst0_O));
Decode2348 Decode2348_inst0(.I(I), .O(Decode2348_inst0_O));
Decode2358 Decode2358_inst0(.I(I), .O(Decode2358_inst0_O));
Decode2368 Decode2368_inst0(.I(I), .O(Decode2368_inst0_O));
Decode2378 Decode2378_inst0(.I(I), .O(Decode2378_inst0_O));
Decode2388 Decode2388_inst0(.I(I), .O(Decode2388_inst0_O));
Decode238 Decode238_inst0(.I(I), .O(Decode238_inst0_O));
Decode2398 Decode2398_inst0(.I(I), .O(Decode2398_inst0_O));
Decode2408 Decode2408_inst0(.I(I), .O(Decode2408_inst0_O));
Decode2418 Decode2418_inst0(.I(I), .O(Decode2418_inst0_O));
Decode2428 Decode2428_inst0(.I(I), .O(Decode2428_inst0_O));
Decode2438 Decode2438_inst0(.I(I), .O(Decode2438_inst0_O));
Decode2448 Decode2448_inst0(.I(I), .O(Decode2448_inst0_O));
Decode2458 Decode2458_inst0(.I(I), .O(Decode2458_inst0_O));
Decode2468 Decode2468_inst0(.I(I), .O(Decode2468_inst0_O));
Decode2478 Decode2478_inst0(.I(I), .O(Decode2478_inst0_O));
Decode2488 Decode2488_inst0(.I(I), .O(Decode2488_inst0_O));
Decode248 Decode248_inst0(.I(I), .O(Decode248_inst0_O));
Decode2498 Decode2498_inst0(.I(I), .O(Decode2498_inst0_O));
Decode2508 Decode2508_inst0(.I(I), .O(Decode2508_inst0_O));
Decode2518 Decode2518_inst0(.I(I), .O(Decode2518_inst0_O));
Decode2528 Decode2528_inst0(.I(I), .O(Decode2528_inst0_O));
Decode2538 Decode2538_inst0(.I(I), .O(Decode2538_inst0_O));
Decode2548 Decode2548_inst0(.I(I), .O(Decode2548_inst0_O));
Decode2558 Decode2558_inst0(.I(I), .O(Decode2558_inst0_O));
Decode258 Decode258_inst0(.I(I), .O(Decode258_inst0_O));
Decode268 Decode268_inst0(.I(I), .O(Decode268_inst0_O));
Decode278 Decode278_inst0(.I(I), .O(Decode278_inst0_O));
Decode288 Decode288_inst0(.I(I), .O(Decode288_inst0_O));
Decode28 Decode28_inst0(.I(I), .O(Decode28_inst0_O));
Decode298 Decode298_inst0(.I(I), .O(Decode298_inst0_O));
Decode308 Decode308_inst0(.I(I), .O(Decode308_inst0_O));
Decode318 Decode318_inst0(.I(I), .O(Decode318_inst0_O));
Decode328 Decode328_inst0(.I(I), .O(Decode328_inst0_O));
Decode338 Decode338_inst0(.I(I), .O(Decode338_inst0_O));
Decode348 Decode348_inst0(.I(I), .O(Decode348_inst0_O));
Decode358 Decode358_inst0(.I(I), .O(Decode358_inst0_O));
Decode368 Decode368_inst0(.I(I), .O(Decode368_inst0_O));
Decode378 Decode378_inst0(.I(I), .O(Decode378_inst0_O));
Decode388 Decode388_inst0(.I(I), .O(Decode388_inst0_O));
Decode38 Decode38_inst0(.I(I), .O(Decode38_inst0_O));
Decode398 Decode398_inst0(.I(I), .O(Decode398_inst0_O));
Decode408 Decode408_inst0(.I(I), .O(Decode408_inst0_O));
Decode418 Decode418_inst0(.I(I), .O(Decode418_inst0_O));
Decode428 Decode428_inst0(.I(I), .O(Decode428_inst0_O));
Decode438 Decode438_inst0(.I(I), .O(Decode438_inst0_O));
Decode448 Decode448_inst0(.I(I), .O(Decode448_inst0_O));
Decode458 Decode458_inst0(.I(I), .O(Decode458_inst0_O));
Decode468 Decode468_inst0(.I(I), .O(Decode468_inst0_O));
Decode478 Decode478_inst0(.I(I), .O(Decode478_inst0_O));
Decode488 Decode488_inst0(.I(I), .O(Decode488_inst0_O));
Decode48 Decode48_inst0(.I(I), .O(Decode48_inst0_O));
Decode498 Decode498_inst0(.I(I), .O(Decode498_inst0_O));
Decode508 Decode508_inst0(.I(I), .O(Decode508_inst0_O));
Decode518 Decode518_inst0(.I(I), .O(Decode518_inst0_O));
Decode528 Decode528_inst0(.I(I), .O(Decode528_inst0_O));
Decode538 Decode538_inst0(.I(I), .O(Decode538_inst0_O));
Decode548 Decode548_inst0(.I(I), .O(Decode548_inst0_O));
Decode558 Decode558_inst0(.I(I), .O(Decode558_inst0_O));
Decode568 Decode568_inst0(.I(I), .O(Decode568_inst0_O));
Decode578 Decode578_inst0(.I(I), .O(Decode578_inst0_O));
Decode588 Decode588_inst0(.I(I), .O(Decode588_inst0_O));
Decode58 Decode58_inst0(.I(I), .O(Decode58_inst0_O));
Decode598 Decode598_inst0(.I(I), .O(Decode598_inst0_O));
Decode608 Decode608_inst0(.I(I), .O(Decode608_inst0_O));
Decode618 Decode618_inst0(.I(I), .O(Decode618_inst0_O));
Decode628 Decode628_inst0(.I(I), .O(Decode628_inst0_O));
Decode638 Decode638_inst0(.I(I), .O(Decode638_inst0_O));
Decode648 Decode648_inst0(.I(I), .O(Decode648_inst0_O));
Decode658 Decode658_inst0(.I(I), .O(Decode658_inst0_O));
Decode668 Decode668_inst0(.I(I), .O(Decode668_inst0_O));
Decode678 Decode678_inst0(.I(I), .O(Decode678_inst0_O));
Decode688 Decode688_inst0(.I(I), .O(Decode688_inst0_O));
Decode68 Decode68_inst0(.I(I), .O(Decode68_inst0_O));
Decode698 Decode698_inst0(.I(I), .O(Decode698_inst0_O));
Decode708 Decode708_inst0(.I(I), .O(Decode708_inst0_O));
Decode718 Decode718_inst0(.I(I), .O(Decode718_inst0_O));
Decode728 Decode728_inst0(.I(I), .O(Decode728_inst0_O));
Decode738 Decode738_inst0(.I(I), .O(Decode738_inst0_O));
Decode748 Decode748_inst0(.I(I), .O(Decode748_inst0_O));
Decode758 Decode758_inst0(.I(I), .O(Decode758_inst0_O));
Decode768 Decode768_inst0(.I(I), .O(Decode768_inst0_O));
Decode778 Decode778_inst0(.I(I), .O(Decode778_inst0_O));
Decode788 Decode788_inst0(.I(I), .O(Decode788_inst0_O));
Decode78 Decode78_inst0(.I(I), .O(Decode78_inst0_O));
Decode798 Decode798_inst0(.I(I), .O(Decode798_inst0_O));
Decode808 Decode808_inst0(.I(I), .O(Decode808_inst0_O));
Decode818 Decode818_inst0(.I(I), .O(Decode818_inst0_O));
Decode828 Decode828_inst0(.I(I), .O(Decode828_inst0_O));
Decode838 Decode838_inst0(.I(I), .O(Decode838_inst0_O));
Decode848 Decode848_inst0(.I(I), .O(Decode848_inst0_O));
Decode858 Decode858_inst0(.I(I), .O(Decode858_inst0_O));
Decode868 Decode868_inst0(.I(I), .O(Decode868_inst0_O));
Decode878 Decode878_inst0(.I(I), .O(Decode878_inst0_O));
Decode888 Decode888_inst0(.I(I), .O(Decode888_inst0_O));
Decode88 Decode88_inst0(.I(I), .O(Decode88_inst0_O));
Decode898 Decode898_inst0(.I(I), .O(Decode898_inst0_O));
Decode908 Decode908_inst0(.I(I), .O(Decode908_inst0_O));
Decode918 Decode918_inst0(.I(I), .O(Decode918_inst0_O));
Decode928 Decode928_inst0(.I(I), .O(Decode928_inst0_O));
Decode938 Decode938_inst0(.I(I), .O(Decode938_inst0_O));
Decode948 Decode948_inst0(.I(I), .O(Decode948_inst0_O));
Decode958 Decode958_inst0(.I(I), .O(Decode958_inst0_O));
Decode968 Decode968_inst0(.I(I), .O(Decode968_inst0_O));
Decode978 Decode978_inst0(.I(I), .O(Decode978_inst0_O));
Decode988 Decode988_inst0(.I(I), .O(Decode988_inst0_O));
Decode98 Decode98_inst0(.I(I), .O(Decode98_inst0_O));
Decode998 Decode998_inst0(.I(I), .O(Decode998_inst0_O));
assign O = {Decode2558_inst0_O,Decode2548_inst0_O,Decode2538_inst0_O,Decode2528_inst0_O,Decode2518_inst0_O,Decode2508_inst0_O,Decode2498_inst0_O,Decode2488_inst0_O,Decode2478_inst0_O,Decode2468_inst0_O,Decode2458_inst0_O,Decode2448_inst0_O,Decode2438_inst0_O,Decode2428_inst0_O,Decode2418_inst0_O,Decode2408_inst0_O,Decode2398_inst0_O,Decode2388_inst0_O,Decode2378_inst0_O,Decode2368_inst0_O,Decode2358_inst0_O,Decode2348_inst0_O,Decode2338_inst0_O,Decode2328_inst0_O,Decode2318_inst0_O,Decode2308_inst0_O,Decode2298_inst0_O,Decode2288_inst0_O,Decode2278_inst0_O,Decode2268_inst0_O,Decode2258_inst0_O,Decode2248_inst0_O,Decode2238_inst0_O,Decode2228_inst0_O,Decode2218_inst0_O,Decode2208_inst0_O,Decode2198_inst0_O,Decode2188_inst0_O,Decode2178_inst0_O,Decode2168_inst0_O,Decode2158_inst0_O,Decode2148_inst0_O,Decode2138_inst0_O,Decode2128_inst0_O,Decode2118_inst0_O,Decode2108_inst0_O,Decode2098_inst0_O,Decode2088_inst0_O,Decode2078_inst0_O,Decode2068_inst0_O,Decode2058_inst0_O,Decode2048_inst0_O,Decode2038_inst0_O,Decode2028_inst0_O,Decode2018_inst0_O,Decode2008_inst0_O,Decode1998_inst0_O,Decode1988_inst0_O,Decode1978_inst0_O,Decode1968_inst0_O,Decode1958_inst0_O,Decode1948_inst0_O,Decode1938_inst0_O,Decode1928_inst0_O,Decode1918_inst0_O,Decode1908_inst0_O,Decode1898_inst0_O,Decode1888_inst0_O,Decode1878_inst0_O,Decode1868_inst0_O,Decode1858_inst0_O,Decode1848_inst0_O,Decode1838_inst0_O,Decode1828_inst0_O,Decode1818_inst0_O,Decode1808_inst0_O,Decode1798_inst0_O,Decode1788_inst0_O,Decode1778_inst0_O,Decode1768_inst0_O,Decode1758_inst0_O,Decode1748_inst0_O,Decode1738_inst0_O,Decode1728_inst0_O,Decode1718_inst0_O,Decode1708_inst0_O,Decode1698_inst0_O,Decode1688_inst0_O,Decode1678_inst0_O,Decode1668_inst0_O,Decode1658_inst0_O,Decode1648_inst0_O,Decode1638_inst0_O,Decode1628_inst0_O,Decode1618_inst0_O,Decode1608_inst0_O,Decode1598_inst0_O,Decode1588_inst0_O,Decode1578_inst0_O,Decode1568_inst0_O,Decode1558_inst0_O,Decode1548_inst0_O,Decode1538_inst0_O,Decode1528_inst0_O,Decode1518_inst0_O,Decode1508_inst0_O,Decode1498_inst0_O,Decode1488_inst0_O,Decode1478_inst0_O,Decode1468_inst0_O,Decode1458_inst0_O,Decode1448_inst0_O,Decode1438_inst0_O,Decode1428_inst0_O,Decode1418_inst0_O,Decode1408_inst0_O,Decode1398_inst0_O,Decode1388_inst0_O,Decode1378_inst0_O,Decode1368_inst0_O,Decode1358_inst0_O,Decode1348_inst0_O,Decode1338_inst0_O,Decode1328_inst0_O,Decode1318_inst0_O,Decode1308_inst0_O,Decode1298_inst0_O,Decode1288_inst0_O,Decode1278_inst0_O,Decode1268_inst0_O,Decode1258_inst0_O,Decode1248_inst0_O,Decode1238_inst0_O,Decode1228_inst0_O,Decode1218_inst0_O,Decode1208_inst0_O,Decode1198_inst0_O,Decode1188_inst0_O,Decode1178_inst0_O,Decode1168_inst0_O,Decode1158_inst0_O,Decode1148_inst0_O,Decode1138_inst0_O,Decode1128_inst0_O,Decode1118_inst0_O,Decode1108_inst0_O,Decode1098_inst0_O,Decode1088_inst0_O,Decode1078_inst0_O,Decode1068_inst0_O,Decode1058_inst0_O,Decode1048_inst0_O,Decode1038_inst0_O,Decode1028_inst0_O,Decode1018_inst0_O,Decode1008_inst0_O,Decode998_inst0_O,Decode988_inst0_O,Decode978_inst0_O,Decode968_inst0_O,Decode958_inst0_O,Decode948_inst0_O,Decode938_inst0_O,Decode928_inst0_O,Decode918_inst0_O,Decode908_inst0_O,Decode898_inst0_O,Decode888_inst0_O,Decode878_inst0_O,Decode868_inst0_O,Decode858_inst0_O,Decode848_inst0_O,Decode838_inst0_O,Decode828_inst0_O,Decode818_inst0_O,Decode808_inst0_O,Decode798_inst0_O,Decode788_inst0_O,Decode778_inst0_O,Decode768_inst0_O,Decode758_inst0_O,Decode748_inst0_O,Decode738_inst0_O,Decode728_inst0_O,Decode718_inst0_O,Decode708_inst0_O,Decode698_inst0_O,Decode688_inst0_O,Decode678_inst0_O,Decode668_inst0_O,Decode658_inst0_O,Decode648_inst0_O,Decode638_inst0_O,Decode628_inst0_O,Decode618_inst0_O,Decode608_inst0_O,Decode598_inst0_O,Decode588_inst0_O,Decode578_inst0_O,Decode568_inst0_O,Decode558_inst0_O,Decode548_inst0_O,Decode538_inst0_O,Decode528_inst0_O,Decode518_inst0_O,Decode508_inst0_O,Decode498_inst0_O,Decode488_inst0_O,Decode478_inst0_O,Decode468_inst0_O,Decode458_inst0_O,Decode448_inst0_O,Decode438_inst0_O,Decode428_inst0_O,Decode418_inst0_O,Decode408_inst0_O,Decode398_inst0_O,Decode388_inst0_O,Decode378_inst0_O,Decode368_inst0_O,Decode358_inst0_O,Decode348_inst0_O,Decode338_inst0_O,Decode328_inst0_O,Decode318_inst0_O,Decode308_inst0_O,Decode298_inst0_O,Decode288_inst0_O,Decode278_inst0_O,Decode268_inst0_O,Decode258_inst0_O,Decode248_inst0_O,Decode238_inst0_O,Decode228_inst0_O,Decode218_inst0_O,Decode208_inst0_O,Decode198_inst0_O,Decode188_inst0_O,Decode178_inst0_O,Decode168_inst0_O,Decode158_inst0_O,Decode148_inst0_O,Decode138_inst0_O,Decode128_inst0_O,Decode118_inst0_O,Decode108_inst0_O,Decode98_inst0_O,Decode88_inst0_O,Decode78_inst0_O,Decode68_inst0_O,Decode58_inst0_O,Decode48_inst0_O,Decode38_inst0_O,Decode28_inst0_O,Decode18_inst0_O,Decode08_inst0_O};
endmodule

