module coreir_eq #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 == in1;
endmodule

module coreir_const #(
    parameter width = 1,
    parameter value = 1
) (
    output [width-1:0] out
);
  assign out = value;
endmodule

module Decode998 (
    input [7:0] I,
    output O
);
wire [7:0] const_99_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h63),
    .width(8)
) const_99_8 (
    .out(const_99_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_99_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode988 (
    input [7:0] I,
    output O
);
wire [7:0] const_98_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h62),
    .width(8)
) const_98_8 (
    .out(const_98_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_98_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode98 (
    input [7:0] I,
    output O
);
wire [7:0] const_9_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_9_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode978 (
    input [7:0] I,
    output O
);
wire [7:0] const_97_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h61),
    .width(8)
) const_97_8 (
    .out(const_97_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_97_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode968 (
    input [7:0] I,
    output O
);
wire [7:0] const_96_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h60),
    .width(8)
) const_96_8 (
    .out(const_96_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_96_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode958 (
    input [7:0] I,
    output O
);
wire [7:0] const_95_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5f),
    .width(8)
) const_95_8 (
    .out(const_95_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_95_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode948 (
    input [7:0] I,
    output O
);
wire [7:0] const_94_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5e),
    .width(8)
) const_94_8 (
    .out(const_94_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_94_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode938 (
    input [7:0] I,
    output O
);
wire [7:0] const_93_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5d),
    .width(8)
) const_93_8 (
    .out(const_93_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_93_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode928 (
    input [7:0] I,
    output O
);
wire [7:0] const_92_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5c),
    .width(8)
) const_92_8 (
    .out(const_92_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_92_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode918 (
    input [7:0] I,
    output O
);
wire [7:0] const_91_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5b),
    .width(8)
) const_91_8 (
    .out(const_91_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_91_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode908 (
    input [7:0] I,
    output O
);
wire [7:0] const_90_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h5a),
    .width(8)
) const_90_8 (
    .out(const_90_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_90_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode898 (
    input [7:0] I,
    output O
);
wire [7:0] const_89_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h59),
    .width(8)
) const_89_8 (
    .out(const_89_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_89_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode888 (
    input [7:0] I,
    output O
);
wire [7:0] const_88_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h58),
    .width(8)
) const_88_8 (
    .out(const_88_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_88_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode88 (
    input [7:0] I,
    output O
);
wire [7:0] const_8_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_8_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode878 (
    input [7:0] I,
    output O
);
wire [7:0] const_87_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h57),
    .width(8)
) const_87_8 (
    .out(const_87_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_87_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode868 (
    input [7:0] I,
    output O
);
wire [7:0] const_86_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h56),
    .width(8)
) const_86_8 (
    .out(const_86_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_86_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode858 (
    input [7:0] I,
    output O
);
wire [7:0] const_85_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h55),
    .width(8)
) const_85_8 (
    .out(const_85_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_85_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode848 (
    input [7:0] I,
    output O
);
wire [7:0] const_84_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h54),
    .width(8)
) const_84_8 (
    .out(const_84_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_84_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode838 (
    input [7:0] I,
    output O
);
wire [7:0] const_83_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h53),
    .width(8)
) const_83_8 (
    .out(const_83_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_83_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode828 (
    input [7:0] I,
    output O
);
wire [7:0] const_82_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h52),
    .width(8)
) const_82_8 (
    .out(const_82_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_82_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode818 (
    input [7:0] I,
    output O
);
wire [7:0] const_81_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h51),
    .width(8)
) const_81_8 (
    .out(const_81_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_81_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode808 (
    input [7:0] I,
    output O
);
wire [7:0] const_80_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h50),
    .width(8)
) const_80_8 (
    .out(const_80_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_80_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode798 (
    input [7:0] I,
    output O
);
wire [7:0] const_79_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4f),
    .width(8)
) const_79_8 (
    .out(const_79_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_79_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode788 (
    input [7:0] I,
    output O
);
wire [7:0] const_78_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4e),
    .width(8)
) const_78_8 (
    .out(const_78_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_78_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode78 (
    input [7:0] I,
    output O
);
wire [7:0] const_7_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_7_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode778 (
    input [7:0] I,
    output O
);
wire [7:0] const_77_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4d),
    .width(8)
) const_77_8 (
    .out(const_77_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_77_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode768 (
    input [7:0] I,
    output O
);
wire [7:0] const_76_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4c),
    .width(8)
) const_76_8 (
    .out(const_76_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_76_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode758 (
    input [7:0] I,
    output O
);
wire [7:0] const_75_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4b),
    .width(8)
) const_75_8 (
    .out(const_75_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_75_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode748 (
    input [7:0] I,
    output O
);
wire [7:0] const_74_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h4a),
    .width(8)
) const_74_8 (
    .out(const_74_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_74_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode738 (
    input [7:0] I,
    output O
);
wire [7:0] const_73_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h49),
    .width(8)
) const_73_8 (
    .out(const_73_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_73_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode728 (
    input [7:0] I,
    output O
);
wire [7:0] const_72_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h48),
    .width(8)
) const_72_8 (
    .out(const_72_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_72_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode718 (
    input [7:0] I,
    output O
);
wire [7:0] const_71_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h47),
    .width(8)
) const_71_8 (
    .out(const_71_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_71_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode708 (
    input [7:0] I,
    output O
);
wire [7:0] const_70_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h46),
    .width(8)
) const_70_8 (
    .out(const_70_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_70_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode698 (
    input [7:0] I,
    output O
);
wire [7:0] const_69_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h45),
    .width(8)
) const_69_8 (
    .out(const_69_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_69_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode688 (
    input [7:0] I,
    output O
);
wire [7:0] const_68_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h44),
    .width(8)
) const_68_8 (
    .out(const_68_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_68_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode68 (
    input [7:0] I,
    output O
);
wire [7:0] const_6_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_6_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode678 (
    input [7:0] I,
    output O
);
wire [7:0] const_67_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h43),
    .width(8)
) const_67_8 (
    .out(const_67_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_67_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode668 (
    input [7:0] I,
    output O
);
wire [7:0] const_66_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h42),
    .width(8)
) const_66_8 (
    .out(const_66_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_66_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode658 (
    input [7:0] I,
    output O
);
wire [7:0] const_65_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h41),
    .width(8)
) const_65_8 (
    .out(const_65_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_65_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode648 (
    input [7:0] I,
    output O
);
wire [7:0] const_64_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h40),
    .width(8)
) const_64_8 (
    .out(const_64_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_64_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode638 (
    input [7:0] I,
    output O
);
wire [7:0] const_63_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3f),
    .width(8)
) const_63_8 (
    .out(const_63_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_63_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode628 (
    input [7:0] I,
    output O
);
wire [7:0] const_62_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3e),
    .width(8)
) const_62_8 (
    .out(const_62_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_62_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode618 (
    input [7:0] I,
    output O
);
wire [7:0] const_61_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3d),
    .width(8)
) const_61_8 (
    .out(const_61_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_61_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode608 (
    input [7:0] I,
    output O
);
wire [7:0] const_60_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3c),
    .width(8)
) const_60_8 (
    .out(const_60_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_60_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode598 (
    input [7:0] I,
    output O
);
wire [7:0] const_59_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3b),
    .width(8)
) const_59_8 (
    .out(const_59_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_59_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode588 (
    input [7:0] I,
    output O
);
wire [7:0] const_58_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h3a),
    .width(8)
) const_58_8 (
    .out(const_58_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_58_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode58 (
    input [7:0] I,
    output O
);
wire [7:0] const_5_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_5_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode578 (
    input [7:0] I,
    output O
);
wire [7:0] const_57_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h39),
    .width(8)
) const_57_8 (
    .out(const_57_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_57_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode568 (
    input [7:0] I,
    output O
);
wire [7:0] const_56_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h38),
    .width(8)
) const_56_8 (
    .out(const_56_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_56_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode558 (
    input [7:0] I,
    output O
);
wire [7:0] const_55_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h37),
    .width(8)
) const_55_8 (
    .out(const_55_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_55_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode548 (
    input [7:0] I,
    output O
);
wire [7:0] const_54_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h36),
    .width(8)
) const_54_8 (
    .out(const_54_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_54_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode538 (
    input [7:0] I,
    output O
);
wire [7:0] const_53_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h35),
    .width(8)
) const_53_8 (
    .out(const_53_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_53_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode528 (
    input [7:0] I,
    output O
);
wire [7:0] const_52_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h34),
    .width(8)
) const_52_8 (
    .out(const_52_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_52_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode518 (
    input [7:0] I,
    output O
);
wire [7:0] const_51_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h33),
    .width(8)
) const_51_8 (
    .out(const_51_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_51_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode508 (
    input [7:0] I,
    output O
);
wire [7:0] const_50_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h32),
    .width(8)
) const_50_8 (
    .out(const_50_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_50_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode498 (
    input [7:0] I,
    output O
);
wire [7:0] const_49_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h31),
    .width(8)
) const_49_8 (
    .out(const_49_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_49_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode488 (
    input [7:0] I,
    output O
);
wire [7:0] const_48_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h30),
    .width(8)
) const_48_8 (
    .out(const_48_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_48_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode48 (
    input [7:0] I,
    output O
);
wire [7:0] const_4_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_4_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode478 (
    input [7:0] I,
    output O
);
wire [7:0] const_47_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2f),
    .width(8)
) const_47_8 (
    .out(const_47_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_47_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode468 (
    input [7:0] I,
    output O
);
wire [7:0] const_46_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2e),
    .width(8)
) const_46_8 (
    .out(const_46_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_46_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode458 (
    input [7:0] I,
    output O
);
wire [7:0] const_45_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2d),
    .width(8)
) const_45_8 (
    .out(const_45_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_45_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode448 (
    input [7:0] I,
    output O
);
wire [7:0] const_44_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2c),
    .width(8)
) const_44_8 (
    .out(const_44_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_44_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode438 (
    input [7:0] I,
    output O
);
wire [7:0] const_43_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2b),
    .width(8)
) const_43_8 (
    .out(const_43_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_43_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode428 (
    input [7:0] I,
    output O
);
wire [7:0] const_42_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h2a),
    .width(8)
) const_42_8 (
    .out(const_42_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_42_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode418 (
    input [7:0] I,
    output O
);
wire [7:0] const_41_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h29),
    .width(8)
) const_41_8 (
    .out(const_41_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_41_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode408 (
    input [7:0] I,
    output O
);
wire [7:0] const_40_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h28),
    .width(8)
) const_40_8 (
    .out(const_40_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_40_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode398 (
    input [7:0] I,
    output O
);
wire [7:0] const_39_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h27),
    .width(8)
) const_39_8 (
    .out(const_39_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_39_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode388 (
    input [7:0] I,
    output O
);
wire [7:0] const_38_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h26),
    .width(8)
) const_38_8 (
    .out(const_38_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_38_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode38 (
    input [7:0] I,
    output O
);
wire [7:0] const_3_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_3_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode378 (
    input [7:0] I,
    output O
);
wire [7:0] const_37_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h25),
    .width(8)
) const_37_8 (
    .out(const_37_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_37_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode368 (
    input [7:0] I,
    output O
);
wire [7:0] const_36_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h24),
    .width(8)
) const_36_8 (
    .out(const_36_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_36_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode358 (
    input [7:0] I,
    output O
);
wire [7:0] const_35_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h23),
    .width(8)
) const_35_8 (
    .out(const_35_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_35_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode348 (
    input [7:0] I,
    output O
);
wire [7:0] const_34_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h22),
    .width(8)
) const_34_8 (
    .out(const_34_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_34_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode338 (
    input [7:0] I,
    output O
);
wire [7:0] const_33_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h21),
    .width(8)
) const_33_8 (
    .out(const_33_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_33_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode328 (
    input [7:0] I,
    output O
);
wire [7:0] const_32_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h20),
    .width(8)
) const_32_8 (
    .out(const_32_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_32_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode318 (
    input [7:0] I,
    output O
);
wire [7:0] const_31_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1f),
    .width(8)
) const_31_8 (
    .out(const_31_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_31_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode308 (
    input [7:0] I,
    output O
);
wire [7:0] const_30_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1e),
    .width(8)
) const_30_8 (
    .out(const_30_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_30_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode298 (
    input [7:0] I,
    output O
);
wire [7:0] const_29_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1d),
    .width(8)
) const_29_8 (
    .out(const_29_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_29_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode288 (
    input [7:0] I,
    output O
);
wire [7:0] const_28_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1c),
    .width(8)
) const_28_8 (
    .out(const_28_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_28_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode28 (
    input [7:0] I,
    output O
);
wire [7:0] const_2_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_2_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode278 (
    input [7:0] I,
    output O
);
wire [7:0] const_27_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1b),
    .width(8)
) const_27_8 (
    .out(const_27_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_27_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode268 (
    input [7:0] I,
    output O
);
wire [7:0] const_26_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h1a),
    .width(8)
) const_26_8 (
    .out(const_26_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_26_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode258 (
    input [7:0] I,
    output O
);
wire [7:0] const_25_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h19),
    .width(8)
) const_25_8 (
    .out(const_25_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_25_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2558 (
    input [7:0] I,
    output O
);
wire [7:0] const_255_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hff),
    .width(8)
) const_255_8 (
    .out(const_255_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_255_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2548 (
    input [7:0] I,
    output O
);
wire [7:0] const_254_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hfe),
    .width(8)
) const_254_8 (
    .out(const_254_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_254_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2538 (
    input [7:0] I,
    output O
);
wire [7:0] const_253_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hfd),
    .width(8)
) const_253_8 (
    .out(const_253_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_253_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2528 (
    input [7:0] I,
    output O
);
wire [7:0] const_252_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hfc),
    .width(8)
) const_252_8 (
    .out(const_252_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_252_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2518 (
    input [7:0] I,
    output O
);
wire [7:0] const_251_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hfb),
    .width(8)
) const_251_8 (
    .out(const_251_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_251_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2508 (
    input [7:0] I,
    output O
);
wire [7:0] const_250_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hfa),
    .width(8)
) const_250_8 (
    .out(const_250_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_250_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2498 (
    input [7:0] I,
    output O
);
wire [7:0] const_249_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf9),
    .width(8)
) const_249_8 (
    .out(const_249_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_249_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2488 (
    input [7:0] I,
    output O
);
wire [7:0] const_248_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf8),
    .width(8)
) const_248_8 (
    .out(const_248_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_248_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode248 (
    input [7:0] I,
    output O
);
wire [7:0] const_24_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h18),
    .width(8)
) const_24_8 (
    .out(const_24_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_24_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2478 (
    input [7:0] I,
    output O
);
wire [7:0] const_247_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf7),
    .width(8)
) const_247_8 (
    .out(const_247_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_247_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2468 (
    input [7:0] I,
    output O
);
wire [7:0] const_246_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf6),
    .width(8)
) const_246_8 (
    .out(const_246_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_246_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2458 (
    input [7:0] I,
    output O
);
wire [7:0] const_245_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf5),
    .width(8)
) const_245_8 (
    .out(const_245_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_245_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2448 (
    input [7:0] I,
    output O
);
wire [7:0] const_244_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf4),
    .width(8)
) const_244_8 (
    .out(const_244_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_244_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2438 (
    input [7:0] I,
    output O
);
wire [7:0] const_243_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf3),
    .width(8)
) const_243_8 (
    .out(const_243_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_243_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2428 (
    input [7:0] I,
    output O
);
wire [7:0] const_242_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf2),
    .width(8)
) const_242_8 (
    .out(const_242_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_242_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2418 (
    input [7:0] I,
    output O
);
wire [7:0] const_241_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf1),
    .width(8)
) const_241_8 (
    .out(const_241_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_241_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2408 (
    input [7:0] I,
    output O
);
wire [7:0] const_240_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hf0),
    .width(8)
) const_240_8 (
    .out(const_240_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_240_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2398 (
    input [7:0] I,
    output O
);
wire [7:0] const_239_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hef),
    .width(8)
) const_239_8 (
    .out(const_239_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_239_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2388 (
    input [7:0] I,
    output O
);
wire [7:0] const_238_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hee),
    .width(8)
) const_238_8 (
    .out(const_238_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_238_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode238 (
    input [7:0] I,
    output O
);
wire [7:0] const_23_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h17),
    .width(8)
) const_23_8 (
    .out(const_23_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_23_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2378 (
    input [7:0] I,
    output O
);
wire [7:0] const_237_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hed),
    .width(8)
) const_237_8 (
    .out(const_237_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_237_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2368 (
    input [7:0] I,
    output O
);
wire [7:0] const_236_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hec),
    .width(8)
) const_236_8 (
    .out(const_236_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_236_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2358 (
    input [7:0] I,
    output O
);
wire [7:0] const_235_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'heb),
    .width(8)
) const_235_8 (
    .out(const_235_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_235_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2348 (
    input [7:0] I,
    output O
);
wire [7:0] const_234_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hea),
    .width(8)
) const_234_8 (
    .out(const_234_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_234_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2338 (
    input [7:0] I,
    output O
);
wire [7:0] const_233_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he9),
    .width(8)
) const_233_8 (
    .out(const_233_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_233_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2328 (
    input [7:0] I,
    output O
);
wire [7:0] const_232_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he8),
    .width(8)
) const_232_8 (
    .out(const_232_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_232_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2318 (
    input [7:0] I,
    output O
);
wire [7:0] const_231_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he7),
    .width(8)
) const_231_8 (
    .out(const_231_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_231_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2308 (
    input [7:0] I,
    output O
);
wire [7:0] const_230_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he6),
    .width(8)
) const_230_8 (
    .out(const_230_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_230_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2298 (
    input [7:0] I,
    output O
);
wire [7:0] const_229_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he5),
    .width(8)
) const_229_8 (
    .out(const_229_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_229_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2288 (
    input [7:0] I,
    output O
);
wire [7:0] const_228_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he4),
    .width(8)
) const_228_8 (
    .out(const_228_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_228_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode228 (
    input [7:0] I,
    output O
);
wire [7:0] const_22_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h16),
    .width(8)
) const_22_8 (
    .out(const_22_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_22_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2278 (
    input [7:0] I,
    output O
);
wire [7:0] const_227_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he3),
    .width(8)
) const_227_8 (
    .out(const_227_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_227_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2268 (
    input [7:0] I,
    output O
);
wire [7:0] const_226_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he2),
    .width(8)
) const_226_8 (
    .out(const_226_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_226_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2258 (
    input [7:0] I,
    output O
);
wire [7:0] const_225_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he1),
    .width(8)
) const_225_8 (
    .out(const_225_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_225_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2248 (
    input [7:0] I,
    output O
);
wire [7:0] const_224_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'he0),
    .width(8)
) const_224_8 (
    .out(const_224_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_224_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2238 (
    input [7:0] I,
    output O
);
wire [7:0] const_223_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hdf),
    .width(8)
) const_223_8 (
    .out(const_223_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_223_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2228 (
    input [7:0] I,
    output O
);
wire [7:0] const_222_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hde),
    .width(8)
) const_222_8 (
    .out(const_222_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_222_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2218 (
    input [7:0] I,
    output O
);
wire [7:0] const_221_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hdd),
    .width(8)
) const_221_8 (
    .out(const_221_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_221_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2208 (
    input [7:0] I,
    output O
);
wire [7:0] const_220_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hdc),
    .width(8)
) const_220_8 (
    .out(const_220_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_220_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2198 (
    input [7:0] I,
    output O
);
wire [7:0] const_219_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hdb),
    .width(8)
) const_219_8 (
    .out(const_219_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_219_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2188 (
    input [7:0] I,
    output O
);
wire [7:0] const_218_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hda),
    .width(8)
) const_218_8 (
    .out(const_218_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_218_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode218 (
    input [7:0] I,
    output O
);
wire [7:0] const_21_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h15),
    .width(8)
) const_21_8 (
    .out(const_21_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_21_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2178 (
    input [7:0] I,
    output O
);
wire [7:0] const_217_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd9),
    .width(8)
) const_217_8 (
    .out(const_217_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_217_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2168 (
    input [7:0] I,
    output O
);
wire [7:0] const_216_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd8),
    .width(8)
) const_216_8 (
    .out(const_216_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_216_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2158 (
    input [7:0] I,
    output O
);
wire [7:0] const_215_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd7),
    .width(8)
) const_215_8 (
    .out(const_215_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_215_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2148 (
    input [7:0] I,
    output O
);
wire [7:0] const_214_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd6),
    .width(8)
) const_214_8 (
    .out(const_214_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_214_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2138 (
    input [7:0] I,
    output O
);
wire [7:0] const_213_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd5),
    .width(8)
) const_213_8 (
    .out(const_213_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_213_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2128 (
    input [7:0] I,
    output O
);
wire [7:0] const_212_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd4),
    .width(8)
) const_212_8 (
    .out(const_212_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_212_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2118 (
    input [7:0] I,
    output O
);
wire [7:0] const_211_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd3),
    .width(8)
) const_211_8 (
    .out(const_211_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_211_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2108 (
    input [7:0] I,
    output O
);
wire [7:0] const_210_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd2),
    .width(8)
) const_210_8 (
    .out(const_210_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_210_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2098 (
    input [7:0] I,
    output O
);
wire [7:0] const_209_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd1),
    .width(8)
) const_209_8 (
    .out(const_209_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_209_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2088 (
    input [7:0] I,
    output O
);
wire [7:0] const_208_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hd0),
    .width(8)
) const_208_8 (
    .out(const_208_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_208_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode208 (
    input [7:0] I,
    output O
);
wire [7:0] const_20_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h14),
    .width(8)
) const_20_8 (
    .out(const_20_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_20_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2078 (
    input [7:0] I,
    output O
);
wire [7:0] const_207_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hcf),
    .width(8)
) const_207_8 (
    .out(const_207_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_207_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2068 (
    input [7:0] I,
    output O
);
wire [7:0] const_206_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hce),
    .width(8)
) const_206_8 (
    .out(const_206_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_206_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2058 (
    input [7:0] I,
    output O
);
wire [7:0] const_205_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hcd),
    .width(8)
) const_205_8 (
    .out(const_205_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_205_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2048 (
    input [7:0] I,
    output O
);
wire [7:0] const_204_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hcc),
    .width(8)
) const_204_8 (
    .out(const_204_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_204_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2038 (
    input [7:0] I,
    output O
);
wire [7:0] const_203_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hcb),
    .width(8)
) const_203_8 (
    .out(const_203_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_203_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2028 (
    input [7:0] I,
    output O
);
wire [7:0] const_202_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hca),
    .width(8)
) const_202_8 (
    .out(const_202_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_202_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2018 (
    input [7:0] I,
    output O
);
wire [7:0] const_201_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc9),
    .width(8)
) const_201_8 (
    .out(const_201_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_201_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode2008 (
    input [7:0] I,
    output O
);
wire [7:0] const_200_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc8),
    .width(8)
) const_200_8 (
    .out(const_200_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_200_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1998 (
    input [7:0] I,
    output O
);
wire [7:0] const_199_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc7),
    .width(8)
) const_199_8 (
    .out(const_199_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_199_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1988 (
    input [7:0] I,
    output O
);
wire [7:0] const_198_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc6),
    .width(8)
) const_198_8 (
    .out(const_198_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_198_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode198 (
    input [7:0] I,
    output O
);
wire [7:0] const_19_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h13),
    .width(8)
) const_19_8 (
    .out(const_19_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_19_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1978 (
    input [7:0] I,
    output O
);
wire [7:0] const_197_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc5),
    .width(8)
) const_197_8 (
    .out(const_197_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_197_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1968 (
    input [7:0] I,
    output O
);
wire [7:0] const_196_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc4),
    .width(8)
) const_196_8 (
    .out(const_196_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_196_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1958 (
    input [7:0] I,
    output O
);
wire [7:0] const_195_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc3),
    .width(8)
) const_195_8 (
    .out(const_195_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_195_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1948 (
    input [7:0] I,
    output O
);
wire [7:0] const_194_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc2),
    .width(8)
) const_194_8 (
    .out(const_194_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_194_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1938 (
    input [7:0] I,
    output O
);
wire [7:0] const_193_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc1),
    .width(8)
) const_193_8 (
    .out(const_193_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_193_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1928 (
    input [7:0] I,
    output O
);
wire [7:0] const_192_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hc0),
    .width(8)
) const_192_8 (
    .out(const_192_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_192_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1918 (
    input [7:0] I,
    output O
);
wire [7:0] const_191_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hbf),
    .width(8)
) const_191_8 (
    .out(const_191_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_191_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1908 (
    input [7:0] I,
    output O
);
wire [7:0] const_190_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hbe),
    .width(8)
) const_190_8 (
    .out(const_190_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_190_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1898 (
    input [7:0] I,
    output O
);
wire [7:0] const_189_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hbd),
    .width(8)
) const_189_8 (
    .out(const_189_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_189_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1888 (
    input [7:0] I,
    output O
);
wire [7:0] const_188_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hbc),
    .width(8)
) const_188_8 (
    .out(const_188_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_188_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode188 (
    input [7:0] I,
    output O
);
wire [7:0] const_18_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h12),
    .width(8)
) const_18_8 (
    .out(const_18_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_18_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1878 (
    input [7:0] I,
    output O
);
wire [7:0] const_187_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hbb),
    .width(8)
) const_187_8 (
    .out(const_187_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_187_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1868 (
    input [7:0] I,
    output O
);
wire [7:0] const_186_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hba),
    .width(8)
) const_186_8 (
    .out(const_186_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_186_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1858 (
    input [7:0] I,
    output O
);
wire [7:0] const_185_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb9),
    .width(8)
) const_185_8 (
    .out(const_185_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_185_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1848 (
    input [7:0] I,
    output O
);
wire [7:0] const_184_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb8),
    .width(8)
) const_184_8 (
    .out(const_184_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_184_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1838 (
    input [7:0] I,
    output O
);
wire [7:0] const_183_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb7),
    .width(8)
) const_183_8 (
    .out(const_183_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_183_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1828 (
    input [7:0] I,
    output O
);
wire [7:0] const_182_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb6),
    .width(8)
) const_182_8 (
    .out(const_182_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_182_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1818 (
    input [7:0] I,
    output O
);
wire [7:0] const_181_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb5),
    .width(8)
) const_181_8 (
    .out(const_181_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_181_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1808 (
    input [7:0] I,
    output O
);
wire [7:0] const_180_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb4),
    .width(8)
) const_180_8 (
    .out(const_180_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_180_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode18 (
    input [7:0] I,
    output O
);
wire [7:0] const_1_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_1_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1798 (
    input [7:0] I,
    output O
);
wire [7:0] const_179_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb3),
    .width(8)
) const_179_8 (
    .out(const_179_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_179_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1788 (
    input [7:0] I,
    output O
);
wire [7:0] const_178_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb2),
    .width(8)
) const_178_8 (
    .out(const_178_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_178_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode178 (
    input [7:0] I,
    output O
);
wire [7:0] const_17_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h11),
    .width(8)
) const_17_8 (
    .out(const_17_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_17_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1778 (
    input [7:0] I,
    output O
);
wire [7:0] const_177_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb1),
    .width(8)
) const_177_8 (
    .out(const_177_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_177_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1768 (
    input [7:0] I,
    output O
);
wire [7:0] const_176_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hb0),
    .width(8)
) const_176_8 (
    .out(const_176_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_176_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1758 (
    input [7:0] I,
    output O
);
wire [7:0] const_175_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'haf),
    .width(8)
) const_175_8 (
    .out(const_175_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_175_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1748 (
    input [7:0] I,
    output O
);
wire [7:0] const_174_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hae),
    .width(8)
) const_174_8 (
    .out(const_174_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_174_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1738 (
    input [7:0] I,
    output O
);
wire [7:0] const_173_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'had),
    .width(8)
) const_173_8 (
    .out(const_173_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_173_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1728 (
    input [7:0] I,
    output O
);
wire [7:0] const_172_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hac),
    .width(8)
) const_172_8 (
    .out(const_172_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_172_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1718 (
    input [7:0] I,
    output O
);
wire [7:0] const_171_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'hab),
    .width(8)
) const_171_8 (
    .out(const_171_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_171_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1708 (
    input [7:0] I,
    output O
);
wire [7:0] const_170_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'haa),
    .width(8)
) const_170_8 (
    .out(const_170_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_170_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1698 (
    input [7:0] I,
    output O
);
wire [7:0] const_169_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha9),
    .width(8)
) const_169_8 (
    .out(const_169_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_169_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1688 (
    input [7:0] I,
    output O
);
wire [7:0] const_168_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha8),
    .width(8)
) const_168_8 (
    .out(const_168_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_168_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode168 (
    input [7:0] I,
    output O
);
wire [7:0] const_16_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_16_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1678 (
    input [7:0] I,
    output O
);
wire [7:0] const_167_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha7),
    .width(8)
) const_167_8 (
    .out(const_167_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_167_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1668 (
    input [7:0] I,
    output O
);
wire [7:0] const_166_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha6),
    .width(8)
) const_166_8 (
    .out(const_166_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_166_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1658 (
    input [7:0] I,
    output O
);
wire [7:0] const_165_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha5),
    .width(8)
) const_165_8 (
    .out(const_165_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_165_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1648 (
    input [7:0] I,
    output O
);
wire [7:0] const_164_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha4),
    .width(8)
) const_164_8 (
    .out(const_164_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_164_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1638 (
    input [7:0] I,
    output O
);
wire [7:0] const_163_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha3),
    .width(8)
) const_163_8 (
    .out(const_163_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_163_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1628 (
    input [7:0] I,
    output O
);
wire [7:0] const_162_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha2),
    .width(8)
) const_162_8 (
    .out(const_162_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_162_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1618 (
    input [7:0] I,
    output O
);
wire [7:0] const_161_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha1),
    .width(8)
) const_161_8 (
    .out(const_161_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_161_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1608 (
    input [7:0] I,
    output O
);
wire [7:0] const_160_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'ha0),
    .width(8)
) const_160_8 (
    .out(const_160_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_160_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1598 (
    input [7:0] I,
    output O
);
wire [7:0] const_159_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9f),
    .width(8)
) const_159_8 (
    .out(const_159_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_159_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1588 (
    input [7:0] I,
    output O
);
wire [7:0] const_158_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9e),
    .width(8)
) const_158_8 (
    .out(const_158_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_158_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode158 (
    input [7:0] I,
    output O
);
wire [7:0] const_15_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_15_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1578 (
    input [7:0] I,
    output O
);
wire [7:0] const_157_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9d),
    .width(8)
) const_157_8 (
    .out(const_157_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_157_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1568 (
    input [7:0] I,
    output O
);
wire [7:0] const_156_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9c),
    .width(8)
) const_156_8 (
    .out(const_156_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_156_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1558 (
    input [7:0] I,
    output O
);
wire [7:0] const_155_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9b),
    .width(8)
) const_155_8 (
    .out(const_155_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_155_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1548 (
    input [7:0] I,
    output O
);
wire [7:0] const_154_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h9a),
    .width(8)
) const_154_8 (
    .out(const_154_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_154_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1538 (
    input [7:0] I,
    output O
);
wire [7:0] const_153_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h99),
    .width(8)
) const_153_8 (
    .out(const_153_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_153_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1528 (
    input [7:0] I,
    output O
);
wire [7:0] const_152_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h98),
    .width(8)
) const_152_8 (
    .out(const_152_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_152_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1518 (
    input [7:0] I,
    output O
);
wire [7:0] const_151_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h97),
    .width(8)
) const_151_8 (
    .out(const_151_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_151_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1508 (
    input [7:0] I,
    output O
);
wire [7:0] const_150_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h96),
    .width(8)
) const_150_8 (
    .out(const_150_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_150_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1498 (
    input [7:0] I,
    output O
);
wire [7:0] const_149_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h95),
    .width(8)
) const_149_8 (
    .out(const_149_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_149_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1488 (
    input [7:0] I,
    output O
);
wire [7:0] const_148_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h94),
    .width(8)
) const_148_8 (
    .out(const_148_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_148_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode148 (
    input [7:0] I,
    output O
);
wire [7:0] const_14_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_14_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1478 (
    input [7:0] I,
    output O
);
wire [7:0] const_147_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h93),
    .width(8)
) const_147_8 (
    .out(const_147_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_147_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1468 (
    input [7:0] I,
    output O
);
wire [7:0] const_146_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h92),
    .width(8)
) const_146_8 (
    .out(const_146_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_146_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1458 (
    input [7:0] I,
    output O
);
wire [7:0] const_145_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h91),
    .width(8)
) const_145_8 (
    .out(const_145_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_145_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1448 (
    input [7:0] I,
    output O
);
wire [7:0] const_144_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h90),
    .width(8)
) const_144_8 (
    .out(const_144_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_144_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1438 (
    input [7:0] I,
    output O
);
wire [7:0] const_143_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8f),
    .width(8)
) const_143_8 (
    .out(const_143_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_143_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1428 (
    input [7:0] I,
    output O
);
wire [7:0] const_142_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8e),
    .width(8)
) const_142_8 (
    .out(const_142_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_142_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1418 (
    input [7:0] I,
    output O
);
wire [7:0] const_141_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8d),
    .width(8)
) const_141_8 (
    .out(const_141_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_141_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1408 (
    input [7:0] I,
    output O
);
wire [7:0] const_140_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8c),
    .width(8)
) const_140_8 (
    .out(const_140_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_140_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1398 (
    input [7:0] I,
    output O
);
wire [7:0] const_139_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8b),
    .width(8)
) const_139_8 (
    .out(const_139_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_139_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1388 (
    input [7:0] I,
    output O
);
wire [7:0] const_138_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h8a),
    .width(8)
) const_138_8 (
    .out(const_138_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_138_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode138 (
    input [7:0] I,
    output O
);
wire [7:0] const_13_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_13_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1378 (
    input [7:0] I,
    output O
);
wire [7:0] const_137_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h89),
    .width(8)
) const_137_8 (
    .out(const_137_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_137_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1368 (
    input [7:0] I,
    output O
);
wire [7:0] const_136_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h88),
    .width(8)
) const_136_8 (
    .out(const_136_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_136_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1358 (
    input [7:0] I,
    output O
);
wire [7:0] const_135_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h87),
    .width(8)
) const_135_8 (
    .out(const_135_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_135_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1348 (
    input [7:0] I,
    output O
);
wire [7:0] const_134_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h86),
    .width(8)
) const_134_8 (
    .out(const_134_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_134_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1338 (
    input [7:0] I,
    output O
);
wire [7:0] const_133_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h85),
    .width(8)
) const_133_8 (
    .out(const_133_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_133_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1328 (
    input [7:0] I,
    output O
);
wire [7:0] const_132_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h84),
    .width(8)
) const_132_8 (
    .out(const_132_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_132_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1318 (
    input [7:0] I,
    output O
);
wire [7:0] const_131_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h83),
    .width(8)
) const_131_8 (
    .out(const_131_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_131_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1308 (
    input [7:0] I,
    output O
);
wire [7:0] const_130_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h82),
    .width(8)
) const_130_8 (
    .out(const_130_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_130_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1298 (
    input [7:0] I,
    output O
);
wire [7:0] const_129_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h81),
    .width(8)
) const_129_8 (
    .out(const_129_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_129_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1288 (
    input [7:0] I,
    output O
);
wire [7:0] const_128_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h80),
    .width(8)
) const_128_8 (
    .out(const_128_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_128_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode128 (
    input [7:0] I,
    output O
);
wire [7:0] const_12_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_12_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1278 (
    input [7:0] I,
    output O
);
wire [7:0] const_127_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7f),
    .width(8)
) const_127_8 (
    .out(const_127_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_127_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1268 (
    input [7:0] I,
    output O
);
wire [7:0] const_126_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7e),
    .width(8)
) const_126_8 (
    .out(const_126_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_126_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1258 (
    input [7:0] I,
    output O
);
wire [7:0] const_125_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7d),
    .width(8)
) const_125_8 (
    .out(const_125_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_125_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1248 (
    input [7:0] I,
    output O
);
wire [7:0] const_124_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7c),
    .width(8)
) const_124_8 (
    .out(const_124_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_124_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1238 (
    input [7:0] I,
    output O
);
wire [7:0] const_123_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7b),
    .width(8)
) const_123_8 (
    .out(const_123_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_123_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1228 (
    input [7:0] I,
    output O
);
wire [7:0] const_122_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h7a),
    .width(8)
) const_122_8 (
    .out(const_122_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_122_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1218 (
    input [7:0] I,
    output O
);
wire [7:0] const_121_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h79),
    .width(8)
) const_121_8 (
    .out(const_121_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_121_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1208 (
    input [7:0] I,
    output O
);
wire [7:0] const_120_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h78),
    .width(8)
) const_120_8 (
    .out(const_120_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_120_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1198 (
    input [7:0] I,
    output O
);
wire [7:0] const_119_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h77),
    .width(8)
) const_119_8 (
    .out(const_119_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_119_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1188 (
    input [7:0] I,
    output O
);
wire [7:0] const_118_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h76),
    .width(8)
) const_118_8 (
    .out(const_118_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_118_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode118 (
    input [7:0] I,
    output O
);
wire [7:0] const_11_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_11_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1178 (
    input [7:0] I,
    output O
);
wire [7:0] const_117_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h75),
    .width(8)
) const_117_8 (
    .out(const_117_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_117_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1168 (
    input [7:0] I,
    output O
);
wire [7:0] const_116_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h74),
    .width(8)
) const_116_8 (
    .out(const_116_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_116_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1158 (
    input [7:0] I,
    output O
);
wire [7:0] const_115_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h73),
    .width(8)
) const_115_8 (
    .out(const_115_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_115_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1148 (
    input [7:0] I,
    output O
);
wire [7:0] const_114_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h72),
    .width(8)
) const_114_8 (
    .out(const_114_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_114_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1138 (
    input [7:0] I,
    output O
);
wire [7:0] const_113_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h71),
    .width(8)
) const_113_8 (
    .out(const_113_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_113_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1128 (
    input [7:0] I,
    output O
);
wire [7:0] const_112_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h70),
    .width(8)
) const_112_8 (
    .out(const_112_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_112_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1118 (
    input [7:0] I,
    output O
);
wire [7:0] const_111_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6f),
    .width(8)
) const_111_8 (
    .out(const_111_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_111_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1108 (
    input [7:0] I,
    output O
);
wire [7:0] const_110_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6e),
    .width(8)
) const_110_8 (
    .out(const_110_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_110_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1098 (
    input [7:0] I,
    output O
);
wire [7:0] const_109_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6d),
    .width(8)
) const_109_8 (
    .out(const_109_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_109_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1088 (
    input [7:0] I,
    output O
);
wire [7:0] const_108_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6c),
    .width(8)
) const_108_8 (
    .out(const_108_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_108_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode108 (
    input [7:0] I,
    output O
);
wire [7:0] const_10_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_10_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1078 (
    input [7:0] I,
    output O
);
wire [7:0] const_107_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6b),
    .width(8)
) const_107_8 (
    .out(const_107_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_107_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1068 (
    input [7:0] I,
    output O
);
wire [7:0] const_106_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h6a),
    .width(8)
) const_106_8 (
    .out(const_106_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_106_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1058 (
    input [7:0] I,
    output O
);
wire [7:0] const_105_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h69),
    .width(8)
) const_105_8 (
    .out(const_105_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_105_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1048 (
    input [7:0] I,
    output O
);
wire [7:0] const_104_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h68),
    .width(8)
) const_104_8 (
    .out(const_104_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_104_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1038 (
    input [7:0] I,
    output O
);
wire [7:0] const_103_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h67),
    .width(8)
) const_103_8 (
    .out(const_103_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_103_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1028 (
    input [7:0] I,
    output O
);
wire [7:0] const_102_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h66),
    .width(8)
) const_102_8 (
    .out(const_102_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_102_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1018 (
    input [7:0] I,
    output O
);
wire [7:0] const_101_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h65),
    .width(8)
) const_101_8 (
    .out(const_101_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_101_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode1008 (
    input [7:0] I,
    output O
);
wire [7:0] const_100_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h64),
    .width(8)
) const_100_8 (
    .out(const_100_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_100_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode08 (
    input [7:0] I,
    output O
);
wire [7:0] const_0_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_0_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decoder8 (
    input [7:0] I,
    output [255:0] O
);
wire Decode08_inst0_O;
wire Decode1008_inst0_O;
wire Decode1018_inst0_O;
wire Decode1028_inst0_O;
wire Decode1038_inst0_O;
wire Decode1048_inst0_O;
wire Decode1058_inst0_O;
wire Decode1068_inst0_O;
wire Decode1078_inst0_O;
wire Decode1088_inst0_O;
wire Decode108_inst0_O;
wire Decode1098_inst0_O;
wire Decode1108_inst0_O;
wire Decode1118_inst0_O;
wire Decode1128_inst0_O;
wire Decode1138_inst0_O;
wire Decode1148_inst0_O;
wire Decode1158_inst0_O;
wire Decode1168_inst0_O;
wire Decode1178_inst0_O;
wire Decode1188_inst0_O;
wire Decode118_inst0_O;
wire Decode1198_inst0_O;
wire Decode1208_inst0_O;
wire Decode1218_inst0_O;
wire Decode1228_inst0_O;
wire Decode1238_inst0_O;
wire Decode1248_inst0_O;
wire Decode1258_inst0_O;
wire Decode1268_inst0_O;
wire Decode1278_inst0_O;
wire Decode1288_inst0_O;
wire Decode128_inst0_O;
wire Decode1298_inst0_O;
wire Decode1308_inst0_O;
wire Decode1318_inst0_O;
wire Decode1328_inst0_O;
wire Decode1338_inst0_O;
wire Decode1348_inst0_O;
wire Decode1358_inst0_O;
wire Decode1368_inst0_O;
wire Decode1378_inst0_O;
wire Decode1388_inst0_O;
wire Decode138_inst0_O;
wire Decode1398_inst0_O;
wire Decode1408_inst0_O;
wire Decode1418_inst0_O;
wire Decode1428_inst0_O;
wire Decode1438_inst0_O;
wire Decode1448_inst0_O;
wire Decode1458_inst0_O;
wire Decode1468_inst0_O;
wire Decode1478_inst0_O;
wire Decode1488_inst0_O;
wire Decode148_inst0_O;
wire Decode1498_inst0_O;
wire Decode1508_inst0_O;
wire Decode1518_inst0_O;
wire Decode1528_inst0_O;
wire Decode1538_inst0_O;
wire Decode1548_inst0_O;
wire Decode1558_inst0_O;
wire Decode1568_inst0_O;
wire Decode1578_inst0_O;
wire Decode1588_inst0_O;
wire Decode158_inst0_O;
wire Decode1598_inst0_O;
wire Decode1608_inst0_O;
wire Decode1618_inst0_O;
wire Decode1628_inst0_O;
wire Decode1638_inst0_O;
wire Decode1648_inst0_O;
wire Decode1658_inst0_O;
wire Decode1668_inst0_O;
wire Decode1678_inst0_O;
wire Decode1688_inst0_O;
wire Decode168_inst0_O;
wire Decode1698_inst0_O;
wire Decode1708_inst0_O;
wire Decode1718_inst0_O;
wire Decode1728_inst0_O;
wire Decode1738_inst0_O;
wire Decode1748_inst0_O;
wire Decode1758_inst0_O;
wire Decode1768_inst0_O;
wire Decode1778_inst0_O;
wire Decode1788_inst0_O;
wire Decode178_inst0_O;
wire Decode1798_inst0_O;
wire Decode1808_inst0_O;
wire Decode1818_inst0_O;
wire Decode1828_inst0_O;
wire Decode1838_inst0_O;
wire Decode1848_inst0_O;
wire Decode1858_inst0_O;
wire Decode1868_inst0_O;
wire Decode1878_inst0_O;
wire Decode1888_inst0_O;
wire Decode188_inst0_O;
wire Decode1898_inst0_O;
wire Decode18_inst0_O;
wire Decode1908_inst0_O;
wire Decode1918_inst0_O;
wire Decode1928_inst0_O;
wire Decode1938_inst0_O;
wire Decode1948_inst0_O;
wire Decode1958_inst0_O;
wire Decode1968_inst0_O;
wire Decode1978_inst0_O;
wire Decode1988_inst0_O;
wire Decode198_inst0_O;
wire Decode1998_inst0_O;
wire Decode2008_inst0_O;
wire Decode2018_inst0_O;
wire Decode2028_inst0_O;
wire Decode2038_inst0_O;
wire Decode2048_inst0_O;
wire Decode2058_inst0_O;
wire Decode2068_inst0_O;
wire Decode2078_inst0_O;
wire Decode2088_inst0_O;
wire Decode208_inst0_O;
wire Decode2098_inst0_O;
wire Decode2108_inst0_O;
wire Decode2118_inst0_O;
wire Decode2128_inst0_O;
wire Decode2138_inst0_O;
wire Decode2148_inst0_O;
wire Decode2158_inst0_O;
wire Decode2168_inst0_O;
wire Decode2178_inst0_O;
wire Decode2188_inst0_O;
wire Decode218_inst0_O;
wire Decode2198_inst0_O;
wire Decode2208_inst0_O;
wire Decode2218_inst0_O;
wire Decode2228_inst0_O;
wire Decode2238_inst0_O;
wire Decode2248_inst0_O;
wire Decode2258_inst0_O;
wire Decode2268_inst0_O;
wire Decode2278_inst0_O;
wire Decode2288_inst0_O;
wire Decode228_inst0_O;
wire Decode2298_inst0_O;
wire Decode2308_inst0_O;
wire Decode2318_inst0_O;
wire Decode2328_inst0_O;
wire Decode2338_inst0_O;
wire Decode2348_inst0_O;
wire Decode2358_inst0_O;
wire Decode2368_inst0_O;
wire Decode2378_inst0_O;
wire Decode2388_inst0_O;
wire Decode238_inst0_O;
wire Decode2398_inst0_O;
wire Decode2408_inst0_O;
wire Decode2418_inst0_O;
wire Decode2428_inst0_O;
wire Decode2438_inst0_O;
wire Decode2448_inst0_O;
wire Decode2458_inst0_O;
wire Decode2468_inst0_O;
wire Decode2478_inst0_O;
wire Decode2488_inst0_O;
wire Decode248_inst0_O;
wire Decode2498_inst0_O;
wire Decode2508_inst0_O;
wire Decode2518_inst0_O;
wire Decode2528_inst0_O;
wire Decode2538_inst0_O;
wire Decode2548_inst0_O;
wire Decode2558_inst0_O;
wire Decode258_inst0_O;
wire Decode268_inst0_O;
wire Decode278_inst0_O;
wire Decode288_inst0_O;
wire Decode28_inst0_O;
wire Decode298_inst0_O;
wire Decode308_inst0_O;
wire Decode318_inst0_O;
wire Decode328_inst0_O;
wire Decode338_inst0_O;
wire Decode348_inst0_O;
wire Decode358_inst0_O;
wire Decode368_inst0_O;
wire Decode378_inst0_O;
wire Decode388_inst0_O;
wire Decode38_inst0_O;
wire Decode398_inst0_O;
wire Decode408_inst0_O;
wire Decode418_inst0_O;
wire Decode428_inst0_O;
wire Decode438_inst0_O;
wire Decode448_inst0_O;
wire Decode458_inst0_O;
wire Decode468_inst0_O;
wire Decode478_inst0_O;
wire Decode488_inst0_O;
wire Decode48_inst0_O;
wire Decode498_inst0_O;
wire Decode508_inst0_O;
wire Decode518_inst0_O;
wire Decode528_inst0_O;
wire Decode538_inst0_O;
wire Decode548_inst0_O;
wire Decode558_inst0_O;
wire Decode568_inst0_O;
wire Decode578_inst0_O;
wire Decode588_inst0_O;
wire Decode58_inst0_O;
wire Decode598_inst0_O;
wire Decode608_inst0_O;
wire Decode618_inst0_O;
wire Decode628_inst0_O;
wire Decode638_inst0_O;
wire Decode648_inst0_O;
wire Decode658_inst0_O;
wire Decode668_inst0_O;
wire Decode678_inst0_O;
wire Decode688_inst0_O;
wire Decode68_inst0_O;
wire Decode698_inst0_O;
wire Decode708_inst0_O;
wire Decode718_inst0_O;
wire Decode728_inst0_O;
wire Decode738_inst0_O;
wire Decode748_inst0_O;
wire Decode758_inst0_O;
wire Decode768_inst0_O;
wire Decode778_inst0_O;
wire Decode788_inst0_O;
wire Decode78_inst0_O;
wire Decode798_inst0_O;
wire Decode808_inst0_O;
wire Decode818_inst0_O;
wire Decode828_inst0_O;
wire Decode838_inst0_O;
wire Decode848_inst0_O;
wire Decode858_inst0_O;
wire Decode868_inst0_O;
wire Decode878_inst0_O;
wire Decode888_inst0_O;
wire Decode88_inst0_O;
wire Decode898_inst0_O;
wire Decode908_inst0_O;
wire Decode918_inst0_O;
wire Decode928_inst0_O;
wire Decode938_inst0_O;
wire Decode948_inst0_O;
wire Decode958_inst0_O;
wire Decode968_inst0_O;
wire Decode978_inst0_O;
wire Decode988_inst0_O;
wire Decode98_inst0_O;
wire Decode998_inst0_O;
Decode08 Decode08_inst0 (
    .I(I),
    .O(Decode08_inst0_O)
);
Decode1008 Decode1008_inst0 (
    .I(I),
    .O(Decode1008_inst0_O)
);
Decode1018 Decode1018_inst0 (
    .I(I),
    .O(Decode1018_inst0_O)
);
Decode1028 Decode1028_inst0 (
    .I(I),
    .O(Decode1028_inst0_O)
);
Decode1038 Decode1038_inst0 (
    .I(I),
    .O(Decode1038_inst0_O)
);
Decode1048 Decode1048_inst0 (
    .I(I),
    .O(Decode1048_inst0_O)
);
Decode1058 Decode1058_inst0 (
    .I(I),
    .O(Decode1058_inst0_O)
);
Decode1068 Decode1068_inst0 (
    .I(I),
    .O(Decode1068_inst0_O)
);
Decode1078 Decode1078_inst0 (
    .I(I),
    .O(Decode1078_inst0_O)
);
Decode1088 Decode1088_inst0 (
    .I(I),
    .O(Decode1088_inst0_O)
);
Decode108 Decode108_inst0 (
    .I(I),
    .O(Decode108_inst0_O)
);
Decode1098 Decode1098_inst0 (
    .I(I),
    .O(Decode1098_inst0_O)
);
Decode1108 Decode1108_inst0 (
    .I(I),
    .O(Decode1108_inst0_O)
);
Decode1118 Decode1118_inst0 (
    .I(I),
    .O(Decode1118_inst0_O)
);
Decode1128 Decode1128_inst0 (
    .I(I),
    .O(Decode1128_inst0_O)
);
Decode1138 Decode1138_inst0 (
    .I(I),
    .O(Decode1138_inst0_O)
);
Decode1148 Decode1148_inst0 (
    .I(I),
    .O(Decode1148_inst0_O)
);
Decode1158 Decode1158_inst0 (
    .I(I),
    .O(Decode1158_inst0_O)
);
Decode1168 Decode1168_inst0 (
    .I(I),
    .O(Decode1168_inst0_O)
);
Decode1178 Decode1178_inst0 (
    .I(I),
    .O(Decode1178_inst0_O)
);
Decode1188 Decode1188_inst0 (
    .I(I),
    .O(Decode1188_inst0_O)
);
Decode118 Decode118_inst0 (
    .I(I),
    .O(Decode118_inst0_O)
);
Decode1198 Decode1198_inst0 (
    .I(I),
    .O(Decode1198_inst0_O)
);
Decode1208 Decode1208_inst0 (
    .I(I),
    .O(Decode1208_inst0_O)
);
Decode1218 Decode1218_inst0 (
    .I(I),
    .O(Decode1218_inst0_O)
);
Decode1228 Decode1228_inst0 (
    .I(I),
    .O(Decode1228_inst0_O)
);
Decode1238 Decode1238_inst0 (
    .I(I),
    .O(Decode1238_inst0_O)
);
Decode1248 Decode1248_inst0 (
    .I(I),
    .O(Decode1248_inst0_O)
);
Decode1258 Decode1258_inst0 (
    .I(I),
    .O(Decode1258_inst0_O)
);
Decode1268 Decode1268_inst0 (
    .I(I),
    .O(Decode1268_inst0_O)
);
Decode1278 Decode1278_inst0 (
    .I(I),
    .O(Decode1278_inst0_O)
);
Decode1288 Decode1288_inst0 (
    .I(I),
    .O(Decode1288_inst0_O)
);
Decode128 Decode128_inst0 (
    .I(I),
    .O(Decode128_inst0_O)
);
Decode1298 Decode1298_inst0 (
    .I(I),
    .O(Decode1298_inst0_O)
);
Decode1308 Decode1308_inst0 (
    .I(I),
    .O(Decode1308_inst0_O)
);
Decode1318 Decode1318_inst0 (
    .I(I),
    .O(Decode1318_inst0_O)
);
Decode1328 Decode1328_inst0 (
    .I(I),
    .O(Decode1328_inst0_O)
);
Decode1338 Decode1338_inst0 (
    .I(I),
    .O(Decode1338_inst0_O)
);
Decode1348 Decode1348_inst0 (
    .I(I),
    .O(Decode1348_inst0_O)
);
Decode1358 Decode1358_inst0 (
    .I(I),
    .O(Decode1358_inst0_O)
);
Decode1368 Decode1368_inst0 (
    .I(I),
    .O(Decode1368_inst0_O)
);
Decode1378 Decode1378_inst0 (
    .I(I),
    .O(Decode1378_inst0_O)
);
Decode1388 Decode1388_inst0 (
    .I(I),
    .O(Decode1388_inst0_O)
);
Decode138 Decode138_inst0 (
    .I(I),
    .O(Decode138_inst0_O)
);
Decode1398 Decode1398_inst0 (
    .I(I),
    .O(Decode1398_inst0_O)
);
Decode1408 Decode1408_inst0 (
    .I(I),
    .O(Decode1408_inst0_O)
);
Decode1418 Decode1418_inst0 (
    .I(I),
    .O(Decode1418_inst0_O)
);
Decode1428 Decode1428_inst0 (
    .I(I),
    .O(Decode1428_inst0_O)
);
Decode1438 Decode1438_inst0 (
    .I(I),
    .O(Decode1438_inst0_O)
);
Decode1448 Decode1448_inst0 (
    .I(I),
    .O(Decode1448_inst0_O)
);
Decode1458 Decode1458_inst0 (
    .I(I),
    .O(Decode1458_inst0_O)
);
Decode1468 Decode1468_inst0 (
    .I(I),
    .O(Decode1468_inst0_O)
);
Decode1478 Decode1478_inst0 (
    .I(I),
    .O(Decode1478_inst0_O)
);
Decode1488 Decode1488_inst0 (
    .I(I),
    .O(Decode1488_inst0_O)
);
Decode148 Decode148_inst0 (
    .I(I),
    .O(Decode148_inst0_O)
);
Decode1498 Decode1498_inst0 (
    .I(I),
    .O(Decode1498_inst0_O)
);
Decode1508 Decode1508_inst0 (
    .I(I),
    .O(Decode1508_inst0_O)
);
Decode1518 Decode1518_inst0 (
    .I(I),
    .O(Decode1518_inst0_O)
);
Decode1528 Decode1528_inst0 (
    .I(I),
    .O(Decode1528_inst0_O)
);
Decode1538 Decode1538_inst0 (
    .I(I),
    .O(Decode1538_inst0_O)
);
Decode1548 Decode1548_inst0 (
    .I(I),
    .O(Decode1548_inst0_O)
);
Decode1558 Decode1558_inst0 (
    .I(I),
    .O(Decode1558_inst0_O)
);
Decode1568 Decode1568_inst0 (
    .I(I),
    .O(Decode1568_inst0_O)
);
Decode1578 Decode1578_inst0 (
    .I(I),
    .O(Decode1578_inst0_O)
);
Decode1588 Decode1588_inst0 (
    .I(I),
    .O(Decode1588_inst0_O)
);
Decode158 Decode158_inst0 (
    .I(I),
    .O(Decode158_inst0_O)
);
Decode1598 Decode1598_inst0 (
    .I(I),
    .O(Decode1598_inst0_O)
);
Decode1608 Decode1608_inst0 (
    .I(I),
    .O(Decode1608_inst0_O)
);
Decode1618 Decode1618_inst0 (
    .I(I),
    .O(Decode1618_inst0_O)
);
Decode1628 Decode1628_inst0 (
    .I(I),
    .O(Decode1628_inst0_O)
);
Decode1638 Decode1638_inst0 (
    .I(I),
    .O(Decode1638_inst0_O)
);
Decode1648 Decode1648_inst0 (
    .I(I),
    .O(Decode1648_inst0_O)
);
Decode1658 Decode1658_inst0 (
    .I(I),
    .O(Decode1658_inst0_O)
);
Decode1668 Decode1668_inst0 (
    .I(I),
    .O(Decode1668_inst0_O)
);
Decode1678 Decode1678_inst0 (
    .I(I),
    .O(Decode1678_inst0_O)
);
Decode1688 Decode1688_inst0 (
    .I(I),
    .O(Decode1688_inst0_O)
);
Decode168 Decode168_inst0 (
    .I(I),
    .O(Decode168_inst0_O)
);
Decode1698 Decode1698_inst0 (
    .I(I),
    .O(Decode1698_inst0_O)
);
Decode1708 Decode1708_inst0 (
    .I(I),
    .O(Decode1708_inst0_O)
);
Decode1718 Decode1718_inst0 (
    .I(I),
    .O(Decode1718_inst0_O)
);
Decode1728 Decode1728_inst0 (
    .I(I),
    .O(Decode1728_inst0_O)
);
Decode1738 Decode1738_inst0 (
    .I(I),
    .O(Decode1738_inst0_O)
);
Decode1748 Decode1748_inst0 (
    .I(I),
    .O(Decode1748_inst0_O)
);
Decode1758 Decode1758_inst0 (
    .I(I),
    .O(Decode1758_inst0_O)
);
Decode1768 Decode1768_inst0 (
    .I(I),
    .O(Decode1768_inst0_O)
);
Decode1778 Decode1778_inst0 (
    .I(I),
    .O(Decode1778_inst0_O)
);
Decode1788 Decode1788_inst0 (
    .I(I),
    .O(Decode1788_inst0_O)
);
Decode178 Decode178_inst0 (
    .I(I),
    .O(Decode178_inst0_O)
);
Decode1798 Decode1798_inst0 (
    .I(I),
    .O(Decode1798_inst0_O)
);
Decode1808 Decode1808_inst0 (
    .I(I),
    .O(Decode1808_inst0_O)
);
Decode1818 Decode1818_inst0 (
    .I(I),
    .O(Decode1818_inst0_O)
);
Decode1828 Decode1828_inst0 (
    .I(I),
    .O(Decode1828_inst0_O)
);
Decode1838 Decode1838_inst0 (
    .I(I),
    .O(Decode1838_inst0_O)
);
Decode1848 Decode1848_inst0 (
    .I(I),
    .O(Decode1848_inst0_O)
);
Decode1858 Decode1858_inst0 (
    .I(I),
    .O(Decode1858_inst0_O)
);
Decode1868 Decode1868_inst0 (
    .I(I),
    .O(Decode1868_inst0_O)
);
Decode1878 Decode1878_inst0 (
    .I(I),
    .O(Decode1878_inst0_O)
);
Decode1888 Decode1888_inst0 (
    .I(I),
    .O(Decode1888_inst0_O)
);
Decode188 Decode188_inst0 (
    .I(I),
    .O(Decode188_inst0_O)
);
Decode1898 Decode1898_inst0 (
    .I(I),
    .O(Decode1898_inst0_O)
);
Decode18 Decode18_inst0 (
    .I(I),
    .O(Decode18_inst0_O)
);
Decode1908 Decode1908_inst0 (
    .I(I),
    .O(Decode1908_inst0_O)
);
Decode1918 Decode1918_inst0 (
    .I(I),
    .O(Decode1918_inst0_O)
);
Decode1928 Decode1928_inst0 (
    .I(I),
    .O(Decode1928_inst0_O)
);
Decode1938 Decode1938_inst0 (
    .I(I),
    .O(Decode1938_inst0_O)
);
Decode1948 Decode1948_inst0 (
    .I(I),
    .O(Decode1948_inst0_O)
);
Decode1958 Decode1958_inst0 (
    .I(I),
    .O(Decode1958_inst0_O)
);
Decode1968 Decode1968_inst0 (
    .I(I),
    .O(Decode1968_inst0_O)
);
Decode1978 Decode1978_inst0 (
    .I(I),
    .O(Decode1978_inst0_O)
);
Decode1988 Decode1988_inst0 (
    .I(I),
    .O(Decode1988_inst0_O)
);
Decode198 Decode198_inst0 (
    .I(I),
    .O(Decode198_inst0_O)
);
Decode1998 Decode1998_inst0 (
    .I(I),
    .O(Decode1998_inst0_O)
);
Decode2008 Decode2008_inst0 (
    .I(I),
    .O(Decode2008_inst0_O)
);
Decode2018 Decode2018_inst0 (
    .I(I),
    .O(Decode2018_inst0_O)
);
Decode2028 Decode2028_inst0 (
    .I(I),
    .O(Decode2028_inst0_O)
);
Decode2038 Decode2038_inst0 (
    .I(I),
    .O(Decode2038_inst0_O)
);
Decode2048 Decode2048_inst0 (
    .I(I),
    .O(Decode2048_inst0_O)
);
Decode2058 Decode2058_inst0 (
    .I(I),
    .O(Decode2058_inst0_O)
);
Decode2068 Decode2068_inst0 (
    .I(I),
    .O(Decode2068_inst0_O)
);
Decode2078 Decode2078_inst0 (
    .I(I),
    .O(Decode2078_inst0_O)
);
Decode2088 Decode2088_inst0 (
    .I(I),
    .O(Decode2088_inst0_O)
);
Decode208 Decode208_inst0 (
    .I(I),
    .O(Decode208_inst0_O)
);
Decode2098 Decode2098_inst0 (
    .I(I),
    .O(Decode2098_inst0_O)
);
Decode2108 Decode2108_inst0 (
    .I(I),
    .O(Decode2108_inst0_O)
);
Decode2118 Decode2118_inst0 (
    .I(I),
    .O(Decode2118_inst0_O)
);
Decode2128 Decode2128_inst0 (
    .I(I),
    .O(Decode2128_inst0_O)
);
Decode2138 Decode2138_inst0 (
    .I(I),
    .O(Decode2138_inst0_O)
);
Decode2148 Decode2148_inst0 (
    .I(I),
    .O(Decode2148_inst0_O)
);
Decode2158 Decode2158_inst0 (
    .I(I),
    .O(Decode2158_inst0_O)
);
Decode2168 Decode2168_inst0 (
    .I(I),
    .O(Decode2168_inst0_O)
);
Decode2178 Decode2178_inst0 (
    .I(I),
    .O(Decode2178_inst0_O)
);
Decode2188 Decode2188_inst0 (
    .I(I),
    .O(Decode2188_inst0_O)
);
Decode218 Decode218_inst0 (
    .I(I),
    .O(Decode218_inst0_O)
);
Decode2198 Decode2198_inst0 (
    .I(I),
    .O(Decode2198_inst0_O)
);
Decode2208 Decode2208_inst0 (
    .I(I),
    .O(Decode2208_inst0_O)
);
Decode2218 Decode2218_inst0 (
    .I(I),
    .O(Decode2218_inst0_O)
);
Decode2228 Decode2228_inst0 (
    .I(I),
    .O(Decode2228_inst0_O)
);
Decode2238 Decode2238_inst0 (
    .I(I),
    .O(Decode2238_inst0_O)
);
Decode2248 Decode2248_inst0 (
    .I(I),
    .O(Decode2248_inst0_O)
);
Decode2258 Decode2258_inst0 (
    .I(I),
    .O(Decode2258_inst0_O)
);
Decode2268 Decode2268_inst0 (
    .I(I),
    .O(Decode2268_inst0_O)
);
Decode2278 Decode2278_inst0 (
    .I(I),
    .O(Decode2278_inst0_O)
);
Decode2288 Decode2288_inst0 (
    .I(I),
    .O(Decode2288_inst0_O)
);
Decode228 Decode228_inst0 (
    .I(I),
    .O(Decode228_inst0_O)
);
Decode2298 Decode2298_inst0 (
    .I(I),
    .O(Decode2298_inst0_O)
);
Decode2308 Decode2308_inst0 (
    .I(I),
    .O(Decode2308_inst0_O)
);
Decode2318 Decode2318_inst0 (
    .I(I),
    .O(Decode2318_inst0_O)
);
Decode2328 Decode2328_inst0 (
    .I(I),
    .O(Decode2328_inst0_O)
);
Decode2338 Decode2338_inst0 (
    .I(I),
    .O(Decode2338_inst0_O)
);
Decode2348 Decode2348_inst0 (
    .I(I),
    .O(Decode2348_inst0_O)
);
Decode2358 Decode2358_inst0 (
    .I(I),
    .O(Decode2358_inst0_O)
);
Decode2368 Decode2368_inst0 (
    .I(I),
    .O(Decode2368_inst0_O)
);
Decode2378 Decode2378_inst0 (
    .I(I),
    .O(Decode2378_inst0_O)
);
Decode2388 Decode2388_inst0 (
    .I(I),
    .O(Decode2388_inst0_O)
);
Decode238 Decode238_inst0 (
    .I(I),
    .O(Decode238_inst0_O)
);
Decode2398 Decode2398_inst0 (
    .I(I),
    .O(Decode2398_inst0_O)
);
Decode2408 Decode2408_inst0 (
    .I(I),
    .O(Decode2408_inst0_O)
);
Decode2418 Decode2418_inst0 (
    .I(I),
    .O(Decode2418_inst0_O)
);
Decode2428 Decode2428_inst0 (
    .I(I),
    .O(Decode2428_inst0_O)
);
Decode2438 Decode2438_inst0 (
    .I(I),
    .O(Decode2438_inst0_O)
);
Decode2448 Decode2448_inst0 (
    .I(I),
    .O(Decode2448_inst0_O)
);
Decode2458 Decode2458_inst0 (
    .I(I),
    .O(Decode2458_inst0_O)
);
Decode2468 Decode2468_inst0 (
    .I(I),
    .O(Decode2468_inst0_O)
);
Decode2478 Decode2478_inst0 (
    .I(I),
    .O(Decode2478_inst0_O)
);
Decode2488 Decode2488_inst0 (
    .I(I),
    .O(Decode2488_inst0_O)
);
Decode248 Decode248_inst0 (
    .I(I),
    .O(Decode248_inst0_O)
);
Decode2498 Decode2498_inst0 (
    .I(I),
    .O(Decode2498_inst0_O)
);
Decode2508 Decode2508_inst0 (
    .I(I),
    .O(Decode2508_inst0_O)
);
Decode2518 Decode2518_inst0 (
    .I(I),
    .O(Decode2518_inst0_O)
);
Decode2528 Decode2528_inst0 (
    .I(I),
    .O(Decode2528_inst0_O)
);
Decode2538 Decode2538_inst0 (
    .I(I),
    .O(Decode2538_inst0_O)
);
Decode2548 Decode2548_inst0 (
    .I(I),
    .O(Decode2548_inst0_O)
);
Decode2558 Decode2558_inst0 (
    .I(I),
    .O(Decode2558_inst0_O)
);
Decode258 Decode258_inst0 (
    .I(I),
    .O(Decode258_inst0_O)
);
Decode268 Decode268_inst0 (
    .I(I),
    .O(Decode268_inst0_O)
);
Decode278 Decode278_inst0 (
    .I(I),
    .O(Decode278_inst0_O)
);
Decode288 Decode288_inst0 (
    .I(I),
    .O(Decode288_inst0_O)
);
Decode28 Decode28_inst0 (
    .I(I),
    .O(Decode28_inst0_O)
);
Decode298 Decode298_inst0 (
    .I(I),
    .O(Decode298_inst0_O)
);
Decode308 Decode308_inst0 (
    .I(I),
    .O(Decode308_inst0_O)
);
Decode318 Decode318_inst0 (
    .I(I),
    .O(Decode318_inst0_O)
);
Decode328 Decode328_inst0 (
    .I(I),
    .O(Decode328_inst0_O)
);
Decode338 Decode338_inst0 (
    .I(I),
    .O(Decode338_inst0_O)
);
Decode348 Decode348_inst0 (
    .I(I),
    .O(Decode348_inst0_O)
);
Decode358 Decode358_inst0 (
    .I(I),
    .O(Decode358_inst0_O)
);
Decode368 Decode368_inst0 (
    .I(I),
    .O(Decode368_inst0_O)
);
Decode378 Decode378_inst0 (
    .I(I),
    .O(Decode378_inst0_O)
);
Decode388 Decode388_inst0 (
    .I(I),
    .O(Decode388_inst0_O)
);
Decode38 Decode38_inst0 (
    .I(I),
    .O(Decode38_inst0_O)
);
Decode398 Decode398_inst0 (
    .I(I),
    .O(Decode398_inst0_O)
);
Decode408 Decode408_inst0 (
    .I(I),
    .O(Decode408_inst0_O)
);
Decode418 Decode418_inst0 (
    .I(I),
    .O(Decode418_inst0_O)
);
Decode428 Decode428_inst0 (
    .I(I),
    .O(Decode428_inst0_O)
);
Decode438 Decode438_inst0 (
    .I(I),
    .O(Decode438_inst0_O)
);
Decode448 Decode448_inst0 (
    .I(I),
    .O(Decode448_inst0_O)
);
Decode458 Decode458_inst0 (
    .I(I),
    .O(Decode458_inst0_O)
);
Decode468 Decode468_inst0 (
    .I(I),
    .O(Decode468_inst0_O)
);
Decode478 Decode478_inst0 (
    .I(I),
    .O(Decode478_inst0_O)
);
Decode488 Decode488_inst0 (
    .I(I),
    .O(Decode488_inst0_O)
);
Decode48 Decode48_inst0 (
    .I(I),
    .O(Decode48_inst0_O)
);
Decode498 Decode498_inst0 (
    .I(I),
    .O(Decode498_inst0_O)
);
Decode508 Decode508_inst0 (
    .I(I),
    .O(Decode508_inst0_O)
);
Decode518 Decode518_inst0 (
    .I(I),
    .O(Decode518_inst0_O)
);
Decode528 Decode528_inst0 (
    .I(I),
    .O(Decode528_inst0_O)
);
Decode538 Decode538_inst0 (
    .I(I),
    .O(Decode538_inst0_O)
);
Decode548 Decode548_inst0 (
    .I(I),
    .O(Decode548_inst0_O)
);
Decode558 Decode558_inst0 (
    .I(I),
    .O(Decode558_inst0_O)
);
Decode568 Decode568_inst0 (
    .I(I),
    .O(Decode568_inst0_O)
);
Decode578 Decode578_inst0 (
    .I(I),
    .O(Decode578_inst0_O)
);
Decode588 Decode588_inst0 (
    .I(I),
    .O(Decode588_inst0_O)
);
Decode58 Decode58_inst0 (
    .I(I),
    .O(Decode58_inst0_O)
);
Decode598 Decode598_inst0 (
    .I(I),
    .O(Decode598_inst0_O)
);
Decode608 Decode608_inst0 (
    .I(I),
    .O(Decode608_inst0_O)
);
Decode618 Decode618_inst0 (
    .I(I),
    .O(Decode618_inst0_O)
);
Decode628 Decode628_inst0 (
    .I(I),
    .O(Decode628_inst0_O)
);
Decode638 Decode638_inst0 (
    .I(I),
    .O(Decode638_inst0_O)
);
Decode648 Decode648_inst0 (
    .I(I),
    .O(Decode648_inst0_O)
);
Decode658 Decode658_inst0 (
    .I(I),
    .O(Decode658_inst0_O)
);
Decode668 Decode668_inst0 (
    .I(I),
    .O(Decode668_inst0_O)
);
Decode678 Decode678_inst0 (
    .I(I),
    .O(Decode678_inst0_O)
);
Decode688 Decode688_inst0 (
    .I(I),
    .O(Decode688_inst0_O)
);
Decode68 Decode68_inst0 (
    .I(I),
    .O(Decode68_inst0_O)
);
Decode698 Decode698_inst0 (
    .I(I),
    .O(Decode698_inst0_O)
);
Decode708 Decode708_inst0 (
    .I(I),
    .O(Decode708_inst0_O)
);
Decode718 Decode718_inst0 (
    .I(I),
    .O(Decode718_inst0_O)
);
Decode728 Decode728_inst0 (
    .I(I),
    .O(Decode728_inst0_O)
);
Decode738 Decode738_inst0 (
    .I(I),
    .O(Decode738_inst0_O)
);
Decode748 Decode748_inst0 (
    .I(I),
    .O(Decode748_inst0_O)
);
Decode758 Decode758_inst0 (
    .I(I),
    .O(Decode758_inst0_O)
);
Decode768 Decode768_inst0 (
    .I(I),
    .O(Decode768_inst0_O)
);
Decode778 Decode778_inst0 (
    .I(I),
    .O(Decode778_inst0_O)
);
Decode788 Decode788_inst0 (
    .I(I),
    .O(Decode788_inst0_O)
);
Decode78 Decode78_inst0 (
    .I(I),
    .O(Decode78_inst0_O)
);
Decode798 Decode798_inst0 (
    .I(I),
    .O(Decode798_inst0_O)
);
Decode808 Decode808_inst0 (
    .I(I),
    .O(Decode808_inst0_O)
);
Decode818 Decode818_inst0 (
    .I(I),
    .O(Decode818_inst0_O)
);
Decode828 Decode828_inst0 (
    .I(I),
    .O(Decode828_inst0_O)
);
Decode838 Decode838_inst0 (
    .I(I),
    .O(Decode838_inst0_O)
);
Decode848 Decode848_inst0 (
    .I(I),
    .O(Decode848_inst0_O)
);
Decode858 Decode858_inst0 (
    .I(I),
    .O(Decode858_inst0_O)
);
Decode868 Decode868_inst0 (
    .I(I),
    .O(Decode868_inst0_O)
);
Decode878 Decode878_inst0 (
    .I(I),
    .O(Decode878_inst0_O)
);
Decode888 Decode888_inst0 (
    .I(I),
    .O(Decode888_inst0_O)
);
Decode88 Decode88_inst0 (
    .I(I),
    .O(Decode88_inst0_O)
);
Decode898 Decode898_inst0 (
    .I(I),
    .O(Decode898_inst0_O)
);
Decode908 Decode908_inst0 (
    .I(I),
    .O(Decode908_inst0_O)
);
Decode918 Decode918_inst0 (
    .I(I),
    .O(Decode918_inst0_O)
);
Decode928 Decode928_inst0 (
    .I(I),
    .O(Decode928_inst0_O)
);
Decode938 Decode938_inst0 (
    .I(I),
    .O(Decode938_inst0_O)
);
Decode948 Decode948_inst0 (
    .I(I),
    .O(Decode948_inst0_O)
);
Decode958 Decode958_inst0 (
    .I(I),
    .O(Decode958_inst0_O)
);
Decode968 Decode968_inst0 (
    .I(I),
    .O(Decode968_inst0_O)
);
Decode978 Decode978_inst0 (
    .I(I),
    .O(Decode978_inst0_O)
);
Decode988 Decode988_inst0 (
    .I(I),
    .O(Decode988_inst0_O)
);
Decode98 Decode98_inst0 (
    .I(I),
    .O(Decode98_inst0_O)
);
Decode998 Decode998_inst0 (
    .I(I),
    .O(Decode998_inst0_O)
);
assign O = {Decode2558_inst0_O,Decode2548_inst0_O,Decode2538_inst0_O,Decode2528_inst0_O,Decode2518_inst0_O,Decode2508_inst0_O,Decode2498_inst0_O,Decode2488_inst0_O,Decode2478_inst0_O,Decode2468_inst0_O,Decode2458_inst0_O,Decode2448_inst0_O,Decode2438_inst0_O,Decode2428_inst0_O,Decode2418_inst0_O,Decode2408_inst0_O,Decode2398_inst0_O,Decode2388_inst0_O,Decode2378_inst0_O,Decode2368_inst0_O,Decode2358_inst0_O,Decode2348_inst0_O,Decode2338_inst0_O,Decode2328_inst0_O,Decode2318_inst0_O,Decode2308_inst0_O,Decode2298_inst0_O,Decode2288_inst0_O,Decode2278_inst0_O,Decode2268_inst0_O,Decode2258_inst0_O,Decode2248_inst0_O,Decode2238_inst0_O,Decode2228_inst0_O,Decode2218_inst0_O,Decode2208_inst0_O,Decode2198_inst0_O,Decode2188_inst0_O,Decode2178_inst0_O,Decode2168_inst0_O,Decode2158_inst0_O,Decode2148_inst0_O,Decode2138_inst0_O,Decode2128_inst0_O,Decode2118_inst0_O,Decode2108_inst0_O,Decode2098_inst0_O,Decode2088_inst0_O,Decode2078_inst0_O,Decode2068_inst0_O,Decode2058_inst0_O,Decode2048_inst0_O,Decode2038_inst0_O,Decode2028_inst0_O,Decode2018_inst0_O,Decode2008_inst0_O,Decode1998_inst0_O,Decode1988_inst0_O,Decode1978_inst0_O,Decode1968_inst0_O,Decode1958_inst0_O,Decode1948_inst0_O,Decode1938_inst0_O,Decode1928_inst0_O,Decode1918_inst0_O,Decode1908_inst0_O,Decode1898_inst0_O,Decode1888_inst0_O,Decode1878_inst0_O,Decode1868_inst0_O,Decode1858_inst0_O,Decode1848_inst0_O,Decode1838_inst0_O,Decode1828_inst0_O,Decode1818_inst0_O,Decode1808_inst0_O,Decode1798_inst0_O,Decode1788_inst0_O,Decode1778_inst0_O,Decode1768_inst0_O,Decode1758_inst0_O,Decode1748_inst0_O,Decode1738_inst0_O,Decode1728_inst0_O,Decode1718_inst0_O,Decode1708_inst0_O,Decode1698_inst0_O,Decode1688_inst0_O,Decode1678_inst0_O,Decode1668_inst0_O,Decode1658_inst0_O,Decode1648_inst0_O,Decode1638_inst0_O,Decode1628_inst0_O,Decode1618_inst0_O,Decode1608_inst0_O,Decode1598_inst0_O,Decode1588_inst0_O,Decode1578_inst0_O,Decode1568_inst0_O,Decode1558_inst0_O,Decode1548_inst0_O,Decode1538_inst0_O,Decode1528_inst0_O,Decode1518_inst0_O,Decode1508_inst0_O,Decode1498_inst0_O,Decode1488_inst0_O,Decode1478_inst0_O,Decode1468_inst0_O,Decode1458_inst0_O,Decode1448_inst0_O,Decode1438_inst0_O,Decode1428_inst0_O,Decode1418_inst0_O,Decode1408_inst0_O,Decode1398_inst0_O,Decode1388_inst0_O,Decode1378_inst0_O,Decode1368_inst0_O,Decode1358_inst0_O,Decode1348_inst0_O,Decode1338_inst0_O,Decode1328_inst0_O,Decode1318_inst0_O,Decode1308_inst0_O,Decode1298_inst0_O,Decode1288_inst0_O,Decode1278_inst0_O,Decode1268_inst0_O,Decode1258_inst0_O,Decode1248_inst0_O,Decode1238_inst0_O,Decode1228_inst0_O,Decode1218_inst0_O,Decode1208_inst0_O,Decode1198_inst0_O,Decode1188_inst0_O,Decode1178_inst0_O,Decode1168_inst0_O,Decode1158_inst0_O,Decode1148_inst0_O,Decode1138_inst0_O,Decode1128_inst0_O,Decode1118_inst0_O,Decode1108_inst0_O,Decode1098_inst0_O,Decode1088_inst0_O,Decode1078_inst0_O,Decode1068_inst0_O,Decode1058_inst0_O,Decode1048_inst0_O,Decode1038_inst0_O,Decode1028_inst0_O,Decode1018_inst0_O,Decode1008_inst0_O,Decode998_inst0_O,Decode988_inst0_O,Decode978_inst0_O,Decode968_inst0_O,Decode958_inst0_O,Decode948_inst0_O,Decode938_inst0_O,Decode928_inst0_O,Decode918_inst0_O,Decode908_inst0_O,Decode898_inst0_O,Decode888_inst0_O,Decode878_inst0_O,Decode868_inst0_O,Decode858_inst0_O,Decode848_inst0_O,Decode838_inst0_O,Decode828_inst0_O,Decode818_inst0_O,Decode808_inst0_O,Decode798_inst0_O,Decode788_inst0_O,Decode778_inst0_O,Decode768_inst0_O,Decode758_inst0_O,Decode748_inst0_O,Decode738_inst0_O,Decode728_inst0_O,Decode718_inst0_O,Decode708_inst0_O,Decode698_inst0_O,Decode688_inst0_O,Decode678_inst0_O,Decode668_inst0_O,Decode658_inst0_O,Decode648_inst0_O,Decode638_inst0_O,Decode628_inst0_O,Decode618_inst0_O,Decode608_inst0_O,Decode598_inst0_O,Decode588_inst0_O,Decode578_inst0_O,Decode568_inst0_O,Decode558_inst0_O,Decode548_inst0_O,Decode538_inst0_O,Decode528_inst0_O,Decode518_inst0_O,Decode508_inst0_O,Decode498_inst0_O,Decode488_inst0_O,Decode478_inst0_O,Decode468_inst0_O,Decode458_inst0_O,Decode448_inst0_O,Decode438_inst0_O,Decode428_inst0_O,Decode418_inst0_O,Decode408_inst0_O,Decode398_inst0_O,Decode388_inst0_O,Decode378_inst0_O,Decode368_inst0_O,Decode358_inst0_O,Decode348_inst0_O,Decode338_inst0_O,Decode328_inst0_O,Decode318_inst0_O,Decode308_inst0_O,Decode298_inst0_O,Decode288_inst0_O,Decode278_inst0_O,Decode268_inst0_O,Decode258_inst0_O,Decode248_inst0_O,Decode238_inst0_O,Decode228_inst0_O,Decode218_inst0_O,Decode208_inst0_O,Decode198_inst0_O,Decode188_inst0_O,Decode178_inst0_O,Decode168_inst0_O,Decode158_inst0_O,Decode148_inst0_O,Decode138_inst0_O,Decode128_inst0_O,Decode118_inst0_O,Decode108_inst0_O,Decode98_inst0_O,Decode88_inst0_O,Decode78_inst0_O,Decode68_inst0_O,Decode58_inst0_O,Decode48_inst0_O,Decode38_inst0_O,Decode28_inst0_O,Decode18_inst0_O,Decode08_inst0_O};
endmodule

