module main (output [7:0] LED, input  CLKIN, input [7:0] SWITCH);
wire [7:0] inst0_DO;
wire [0:0] inst0_DOP;
RAMB16_S9 #(.INIT_39(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_2A(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_2B(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_2C(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_2D(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_2E(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_2F(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_0B(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_0C(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_0A(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_0F(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_0D(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_0E(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.WRITE_MODE("WRITE_FIRST"),
.INIT_15(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_14(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_17(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_16(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_11(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_10(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_13(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_12(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_19(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_18(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT(9'h000),
.INIT_38(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_32(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_37(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_36(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_35(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_34(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_05(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.SRVAL(9'h000),
.INIT_3C(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_3B(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_3A(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_01(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_3F(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_3E(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_3D(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_1E(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_33(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_1F(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_1A(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_1C(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_1B(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_31(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_02(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_03(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_00(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_30(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_06(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_07(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_04(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_1D(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INITP_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_08(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_09(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INITP_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_28(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_29(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INITP_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_23(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0),
.INIT_20(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_21(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_22(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INITP_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
.INIT_24(256'h3E3C3A38363432302E2C2A28262422201E1C1A18161412100E0C0A0806040200),
.INIT_25(256'h7E7C7A78767472706E6C6A68666462605E5C5A58565452504E4C4A4846444240),
.INIT_26(256'hBEBCBAB8B6B4B2B0AEACAAA8A6A4A2A09E9C9A98969492908E8C8A8886848280),
.INIT_27(256'hFEFCFAF8F6F4F2F0EEECEAE8E6E4E2E0DEDCDAD8D6D4D2D0CECCCAC8C6C4C2C0)) inst0 (.DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .DIP({1'b0}), .DO(inst0_DO), .DOP(inst0_DOP), .ADDR({1'b0,1'b0,1'b0,SWITCH[7],SWITCH[6],SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .CLK(CLKIN), .EN(1'b1), .SSR(1'b0), .WE(1'b0));
assign LED = {inst0_DOP[0],inst0_DO[7],inst0_DO[6],inst0_DO[5],inst0_DO[4],inst0_DO[3],inst0_DO[2],inst0_DO[1]};
endmodule

