module Adders24_2_2_cin1_cout1 (input [23:0] I0, output [23:0] O, input  CIN, output  COUT);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
wire  inst64_O;
wire  inst65_O;
wire  inst66_O;
wire  inst67_O;
wire  inst68_O;
wire  inst69_O;
wire  inst70_O;
wire  inst71_O;
LUT1 #(.INIT(2'h2)) inst0 (.I0(I0[0]), .O(inst0_O));
MUXCY inst1 (.DI(I0[0]), .CI(CIN), .S(inst0_O), .O(inst1_O));
XORCY inst2 (.LI(inst0_O), .CI(CIN), .O(inst2_O));
LUT1 #(.INIT(2'h2)) inst3 (.I0(I0[1]), .O(inst3_O));
MUXCY inst4 (.DI(I0[1]), .CI(inst1_O), .S(inst3_O), .O(inst4_O));
XORCY inst5 (.LI(inst3_O), .CI(inst1_O), .O(inst5_O));
LUT1 #(.INIT(2'h2)) inst6 (.I0(I0[2]), .O(inst6_O));
MUXCY inst7 (.DI(I0[2]), .CI(inst4_O), .S(inst6_O), .O(inst7_O));
XORCY inst8 (.LI(inst6_O), .CI(inst4_O), .O(inst8_O));
LUT1 #(.INIT(2'h2)) inst9 (.I0(I0[3]), .O(inst9_O));
MUXCY inst10 (.DI(I0[3]), .CI(inst7_O), .S(inst9_O), .O(inst10_O));
XORCY inst11 (.LI(inst9_O), .CI(inst7_O), .O(inst11_O));
LUT1 #(.INIT(2'h2)) inst12 (.I0(I0[4]), .O(inst12_O));
MUXCY inst13 (.DI(I0[4]), .CI(inst10_O), .S(inst12_O), .O(inst13_O));
XORCY inst14 (.LI(inst12_O), .CI(inst10_O), .O(inst14_O));
LUT1 #(.INIT(2'h2)) inst15 (.I0(I0[5]), .O(inst15_O));
MUXCY inst16 (.DI(I0[5]), .CI(inst13_O), .S(inst15_O), .O(inst16_O));
XORCY inst17 (.LI(inst15_O), .CI(inst13_O), .O(inst17_O));
LUT1 #(.INIT(2'h2)) inst18 (.I0(I0[6]), .O(inst18_O));
MUXCY inst19 (.DI(I0[6]), .CI(inst16_O), .S(inst18_O), .O(inst19_O));
XORCY inst20 (.LI(inst18_O), .CI(inst16_O), .O(inst20_O));
LUT1 #(.INIT(2'h2)) inst21 (.I0(I0[7]), .O(inst21_O));
MUXCY inst22 (.DI(I0[7]), .CI(inst19_O), .S(inst21_O), .O(inst22_O));
XORCY inst23 (.LI(inst21_O), .CI(inst19_O), .O(inst23_O));
LUT1 #(.INIT(2'h2)) inst24 (.I0(I0[8]), .O(inst24_O));
MUXCY inst25 (.DI(I0[8]), .CI(inst22_O), .S(inst24_O), .O(inst25_O));
XORCY inst26 (.LI(inst24_O), .CI(inst22_O), .O(inst26_O));
LUT1 #(.INIT(2'h2)) inst27 (.I0(I0[9]), .O(inst27_O));
MUXCY inst28 (.DI(I0[9]), .CI(inst25_O), .S(inst27_O), .O(inst28_O));
XORCY inst29 (.LI(inst27_O), .CI(inst25_O), .O(inst29_O));
LUT1 #(.INIT(2'h2)) inst30 (.I0(I0[10]), .O(inst30_O));
MUXCY inst31 (.DI(I0[10]), .CI(inst28_O), .S(inst30_O), .O(inst31_O));
XORCY inst32 (.LI(inst30_O), .CI(inst28_O), .O(inst32_O));
LUT1 #(.INIT(2'h2)) inst33 (.I0(I0[11]), .O(inst33_O));
MUXCY inst34 (.DI(I0[11]), .CI(inst31_O), .S(inst33_O), .O(inst34_O));
XORCY inst35 (.LI(inst33_O), .CI(inst31_O), .O(inst35_O));
LUT1 #(.INIT(2'h2)) inst36 (.I0(I0[12]), .O(inst36_O));
MUXCY inst37 (.DI(I0[12]), .CI(inst34_O), .S(inst36_O), .O(inst37_O));
XORCY inst38 (.LI(inst36_O), .CI(inst34_O), .O(inst38_O));
LUT1 #(.INIT(2'h2)) inst39 (.I0(I0[13]), .O(inst39_O));
MUXCY inst40 (.DI(I0[13]), .CI(inst37_O), .S(inst39_O), .O(inst40_O));
XORCY inst41 (.LI(inst39_O), .CI(inst37_O), .O(inst41_O));
LUT1 #(.INIT(2'h2)) inst42 (.I0(I0[14]), .O(inst42_O));
MUXCY inst43 (.DI(I0[14]), .CI(inst40_O), .S(inst42_O), .O(inst43_O));
XORCY inst44 (.LI(inst42_O), .CI(inst40_O), .O(inst44_O));
LUT1 #(.INIT(2'h2)) inst45 (.I0(I0[15]), .O(inst45_O));
MUXCY inst46 (.DI(I0[15]), .CI(inst43_O), .S(inst45_O), .O(inst46_O));
XORCY inst47 (.LI(inst45_O), .CI(inst43_O), .O(inst47_O));
LUT1 #(.INIT(2'h2)) inst48 (.I0(I0[16]), .O(inst48_O));
MUXCY inst49 (.DI(I0[16]), .CI(inst46_O), .S(inst48_O), .O(inst49_O));
XORCY inst50 (.LI(inst48_O), .CI(inst46_O), .O(inst50_O));
LUT1 #(.INIT(2'h2)) inst51 (.I0(I0[17]), .O(inst51_O));
MUXCY inst52 (.DI(I0[17]), .CI(inst49_O), .S(inst51_O), .O(inst52_O));
XORCY inst53 (.LI(inst51_O), .CI(inst49_O), .O(inst53_O));
LUT1 #(.INIT(2'h2)) inst54 (.I0(I0[18]), .O(inst54_O));
MUXCY inst55 (.DI(I0[18]), .CI(inst52_O), .S(inst54_O), .O(inst55_O));
XORCY inst56 (.LI(inst54_O), .CI(inst52_O), .O(inst56_O));
LUT1 #(.INIT(2'h2)) inst57 (.I0(I0[19]), .O(inst57_O));
MUXCY inst58 (.DI(I0[19]), .CI(inst55_O), .S(inst57_O), .O(inst58_O));
XORCY inst59 (.LI(inst57_O), .CI(inst55_O), .O(inst59_O));
LUT1 #(.INIT(2'h2)) inst60 (.I0(I0[20]), .O(inst60_O));
MUXCY inst61 (.DI(I0[20]), .CI(inst58_O), .S(inst60_O), .O(inst61_O));
XORCY inst62 (.LI(inst60_O), .CI(inst58_O), .O(inst62_O));
LUT1 #(.INIT(2'h2)) inst63 (.I0(I0[21]), .O(inst63_O));
MUXCY inst64 (.DI(I0[21]), .CI(inst61_O), .S(inst63_O), .O(inst64_O));
XORCY inst65 (.LI(inst63_O), .CI(inst61_O), .O(inst65_O));
LUT1 #(.INIT(2'h2)) inst66 (.I0(I0[22]), .O(inst66_O));
MUXCY inst67 (.DI(I0[22]), .CI(inst64_O), .S(inst66_O), .O(inst67_O));
XORCY inst68 (.LI(inst66_O), .CI(inst64_O), .O(inst68_O));
LUT1 #(.INIT(2'h2)) inst69 (.I0(I0[23]), .O(inst69_O));
MUXCY inst70 (.DI(I0[23]), .CI(inst67_O), .S(inst69_O), .O(inst70_O));
XORCY inst71 (.LI(inst69_O), .CI(inst67_O), .O(inst71_O));
assign O = {inst71_O,inst68_O,inst65_O,inst62_O,inst59_O,inst56_O,inst53_O,inst50_O,inst47_O,inst44_O,inst41_O,inst38_O,inst35_O,inst32_O,inst29_O,inst26_O,inst23_O,inst20_O,inst17_O,inst14_O,inst11_O,inst8_O,inst5_O,inst2_O};
assign COUT = inst70_O;
endmodule

module Register24 (input [23:0] I, output [23:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
wire  inst16_Q;
wire  inst17_Q;
wire  inst18_Q;
wire  inst19_Q;
wire  inst20_Q;
wire  inst21_Q;
wire  inst22_Q;
wire  inst23_Q;
FDRSE #(.INIT(1'h0)) inst0 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[0]), .Q(inst0_Q));
FDRSE #(.INIT(1'h0)) inst1 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[1]), .Q(inst1_Q));
FDRSE #(.INIT(1'h0)) inst2 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[2]), .Q(inst2_Q));
FDRSE #(.INIT(1'h0)) inst3 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[3]), .Q(inst3_Q));
FDRSE #(.INIT(1'h0)) inst4 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[4]), .Q(inst4_Q));
FDRSE #(.INIT(1'h0)) inst5 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[5]), .Q(inst5_Q));
FDRSE #(.INIT(1'h0)) inst6 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[6]), .Q(inst6_Q));
FDRSE #(.INIT(1'h0)) inst7 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[7]), .Q(inst7_Q));
FDRSE #(.INIT(1'h0)) inst8 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[8]), .Q(inst8_Q));
FDRSE #(.INIT(1'h0)) inst9 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[9]), .Q(inst9_Q));
FDRSE #(.INIT(1'h0)) inst10 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[10]), .Q(inst10_Q));
FDRSE #(.INIT(1'h0)) inst11 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[11]), .Q(inst11_Q));
FDRSE #(.INIT(1'h0)) inst12 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[12]), .Q(inst12_Q));
FDRSE #(.INIT(1'h0)) inst13 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[13]), .Q(inst13_Q));
FDRSE #(.INIT(1'h0)) inst14 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[14]), .Q(inst14_Q));
FDRSE #(.INIT(1'h0)) inst15 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[15]), .Q(inst15_Q));
FDRSE #(.INIT(1'h0)) inst16 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[16]), .Q(inst16_Q));
FDRSE #(.INIT(1'h0)) inst17 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[17]), .Q(inst17_Q));
FDRSE #(.INIT(1'h0)) inst18 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[18]), .Q(inst18_Q));
FDRSE #(.INIT(1'h0)) inst19 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[19]), .Q(inst19_Q));
FDRSE #(.INIT(1'h0)) inst20 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[20]), .Q(inst20_Q));
FDRSE #(.INIT(1'h0)) inst21 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[21]), .Q(inst21_Q));
FDRSE #(.INIT(1'h0)) inst22 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[22]), .Q(inst22_Q));
FDRSE #(.INIT(1'h0)) inst23 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[23]), .Q(inst23_Q));
assign O = {inst23_Q,inst22_Q,inst21_Q,inst20_Q,inst19_Q,inst18_Q,inst17_Q,inst16_Q,inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter24_AAAA_AAAA (output [23:0] O, output  COUT, input  CLK);
wire [23:0] inst0_O;
wire  inst0_COUT;
wire [23:0] inst1_O;
Adders24_2_2_cin1_cout1 inst0 (.I0(inst1_O), .O(inst0_O), .CIN(1'b1), .COUT(inst0_COUT));
Register24 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Register4CE_1 (input [3:0] I, output [3:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
FDRSE #(.INIT(1'h1)) inst0 (.C(CLK), .CE(CE), .R(1'b0), .S(1'b0), .D(I[0]), .Q(inst0_Q));
FDRSE #(.INIT(1'h0)) inst1 (.C(CLK), .CE(CE), .R(1'b0), .S(1'b0), .D(I[1]), .Q(inst1_Q));
FDRSE #(.INIT(1'h0)) inst2 (.C(CLK), .CE(CE), .R(1'b0), .S(1'b0), .D(I[2]), .Q(inst2_Q));
FDRSE #(.INIT(1'h0)) inst3 (.C(CLK), .CE(CE), .R(1'b0), .S(1'b0), .D(I[3]), .Q(inst3_Q));
assign O = {inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module PISO4CE_1 (input  SI, input [3:0] PI, input  LOAD, output  O, input  CLK, input  CE);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire [3:0] inst4_O;
LUT3 #(.INIT(8'hCA)) inst0 (.I0(SI), .I1(PI[0]), .I2(LOAD), .O(inst0_O));
LUT3 #(.INIT(8'hCA)) inst1 (.I0(inst4_O[0]), .I1(PI[1]), .I2(LOAD), .O(inst1_O));
LUT3 #(.INIT(8'hCA)) inst2 (.I0(inst4_O[1]), .I1(PI[2]), .I2(LOAD), .O(inst2_O));
LUT3 #(.INIT(8'hCA)) inst3 (.I0(inst4_O[2]), .I1(PI[3]), .I2(LOAD), .O(inst3_O));
Register4CE_1 inst4 (.I({inst3_O,inst2_O,inst1_O,inst0_O}), .O(inst4_O), .CLK(CLK), .CE(CE));
assign O = inst4_O[3];
endmodule

module main (output [0:0] LED, input  CLKIN, input [5:0] SWITCH);
wire [23:0] inst0_O;
wire  inst0_COUT;
wire  inst1_O;
Counter24_AAAA_AAAA inst0 (.O(inst0_O), .COUT(inst0_COUT), .CLK(CLKIN));
PISO4CE_1 inst1 (.SI(SWITCH[0]), .PI({SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1]}), .LOAD(SWITCH[5]), .O(inst1_O), .CLK(CLKIN), .CE(inst0_COUT));
assign LED = {inst1_O};
endmodule

