module main (input  I, output  O);
wire  inst0_0;
not inst0 (inst0_0, I);
assign O = inst0_0;
endmodule

