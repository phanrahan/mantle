module Decode8 (input [7:0] I, output  O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
LUT4 #(.INIT(16'h0001)) inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst0_O));
LUT4 #(.INIT(16'h0000)) inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst1_O));
MUXF5 inst2 (.I0(inst0_O), .I1(inst1_O), .S(I[4]), .O(inst2_O));
LUT4 #(.INIT(16'h0000)) inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst3_O));
LUT4 #(.INIT(16'h0000)) inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst4_O));
MUXF5 inst5 (.I0(inst3_O), .I1(inst4_O), .S(I[4]), .O(inst5_O));
MUXF6 inst6 (.I0(inst2_O), .I1(inst5_O), .S(I[5]), .O(inst6_O));
LUT4 #(.INIT(16'h0000)) inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst7_O));
LUT4 #(.INIT(16'h0000)) inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst8_O));
MUXF5 inst9 (.I0(inst7_O), .I1(inst8_O), .S(I[4]), .O(inst9_O));
LUT4 #(.INIT(16'h0000)) inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst10_O));
LUT4 #(.INIT(16'h0000)) inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst11_O));
MUXF5 inst12 (.I0(inst10_O), .I1(inst11_O), .S(I[4]), .O(inst12_O));
MUXF6 inst13 (.I0(inst9_O), .I1(inst12_O), .S(I[5]), .O(inst13_O));
MUXF7 inst14 (.I0(inst6_O), .I1(inst13_O), .S(I[6]), .O(inst14_O));
LUT4 #(.INIT(16'h0000)) inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst15_O));
LUT4 #(.INIT(16'h0000)) inst16 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst16_O));
MUXF5 inst17 (.I0(inst15_O), .I1(inst16_O), .S(I[4]), .O(inst17_O));
LUT4 #(.INIT(16'h0000)) inst18 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst18_O));
LUT4 #(.INIT(16'h0000)) inst19 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst19_O));
MUXF5 inst20 (.I0(inst18_O), .I1(inst19_O), .S(I[4]), .O(inst20_O));
MUXF6 inst21 (.I0(inst17_O), .I1(inst20_O), .S(I[5]), .O(inst21_O));
LUT4 #(.INIT(16'h0000)) inst22 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst22_O));
LUT4 #(.INIT(16'h0000)) inst23 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst23_O));
MUXF5 inst24 (.I0(inst22_O), .I1(inst23_O), .S(I[4]), .O(inst24_O));
LUT4 #(.INIT(16'h0000)) inst25 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst25_O));
LUT4 #(.INIT(16'h0000)) inst26 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst26_O));
MUXF5 inst27 (.I0(inst25_O), .I1(inst26_O), .S(I[4]), .O(inst27_O));
MUXF6 inst28 (.I0(inst24_O), .I1(inst27_O), .S(I[5]), .O(inst28_O));
MUXF7 inst29 (.I0(inst21_O), .I1(inst28_O), .S(I[6]), .O(inst29_O));
MUXF8 inst30 (.I0(inst14_O), .I1(inst29_O), .S(I[7]), .O(inst30_O));
assign O = inst30_O;
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
wire  inst64_O;
wire  inst65_O;
wire  inst66_O;
wire  inst67_O;
wire  inst68_O;
wire  inst69_O;
wire  inst70_O;
wire  inst71_O;
wire  inst72_O;
wire  inst73_O;
wire  inst74_O;
wire  inst75_O;
wire  inst76_O;
wire  inst77_O;
wire  inst78_O;
wire  inst79_O;
wire  inst80_O;
wire  inst81_O;
wire  inst82_O;
wire  inst83_O;
wire  inst84_O;
wire  inst85_O;
wire  inst86_O;
wire  inst87_O;
wire  inst88_O;
wire  inst89_O;
wire  inst90_O;
wire  inst91_O;
wire  inst92_O;
wire  inst93_O;
wire  inst94_O;
wire  inst95_O;
wire  inst96_O;
wire  inst97_O;
wire  inst98_O;
wire  inst99_O;
wire  inst100_O;
wire  inst101_O;
wire  inst102_O;
wire  inst103_O;
wire  inst104_O;
wire  inst105_O;
wire  inst106_O;
wire  inst107_O;
wire  inst108_O;
wire  inst109_O;
wire  inst110_O;
wire  inst111_O;
wire  inst112_O;
wire  inst113_O;
wire  inst114_O;
wire  inst115_O;
wire  inst116_O;
wire  inst117_O;
wire  inst118_O;
wire  inst119_O;
wire  inst120_O;
wire  inst121_O;
wire  inst122_O;
wire  inst123_O;
wire  inst124_O;
wire  inst125_O;
wire  inst126_O;
wire  inst127_O;
wire  inst128_O;
wire  inst129_O;
wire  inst130_O;
wire  inst131_O;
wire  inst132_O;
wire  inst133_O;
wire  inst134_O;
wire  inst135_O;
wire  inst136_O;
wire  inst137_O;
wire  inst138_O;
wire  inst139_O;
wire  inst140_O;
wire  inst141_O;
wire  inst142_O;
wire  inst143_O;
wire  inst144_O;
wire  inst145_O;
wire  inst146_O;
wire  inst147_O;
wire  inst148_O;
wire  inst149_O;
wire  inst150_O;
wire  inst151_O;
wire  inst152_O;
wire  inst153_O;
wire  inst154_O;
wire  inst155_O;
wire  inst156_O;
wire  inst157_O;
wire  inst158_O;
wire  inst159_O;
wire  inst160_O;
wire  inst161_O;
wire  inst162_O;
wire  inst163_O;
wire  inst164_O;
wire  inst165_O;
wire  inst166_O;
wire  inst167_O;
wire  inst168_O;
wire  inst169_O;
wire  inst170_O;
wire  inst171_O;
wire  inst172_O;
wire  inst173_O;
wire  inst174_O;
wire  inst175_O;
wire  inst176_O;
wire  inst177_O;
wire  inst178_O;
wire  inst179_O;
wire  inst180_O;
wire  inst181_O;
wire  inst182_O;
wire  inst183_O;
wire  inst184_O;
wire  inst185_O;
wire  inst186_O;
wire  inst187_O;
wire  inst188_O;
wire  inst189_O;
wire  inst190_O;
wire  inst191_O;
wire  inst192_O;
wire  inst193_O;
wire  inst194_O;
wire  inst195_O;
wire  inst196_O;
wire  inst197_O;
wire  inst198_O;
wire  inst199_O;
wire  inst200_O;
wire  inst201_O;
wire  inst202_O;
wire  inst203_O;
wire  inst204_O;
wire  inst205_O;
wire  inst206_O;
wire  inst207_O;
wire  inst208_O;
wire  inst209_O;
wire  inst210_O;
wire  inst211_O;
wire  inst212_O;
wire  inst213_O;
wire  inst214_O;
wire  inst215_O;
wire  inst216_O;
wire  inst217_O;
wire  inst218_O;
wire  inst219_O;
wire  inst220_O;
wire  inst221_O;
wire  inst222_O;
wire  inst223_O;
wire  inst224_O;
wire  inst225_O;
wire  inst226_O;
wire  inst227_O;
wire  inst228_O;
wire  inst229_O;
wire  inst230_O;
wire  inst231_O;
wire  inst232_O;
wire  inst233_O;
wire  inst234_O;
wire  inst235_O;
wire  inst236_O;
wire  inst237_O;
wire  inst238_O;
wire  inst239_O;
wire  inst240_O;
wire  inst241_O;
wire  inst242_O;
wire  inst243_O;
wire  inst244_O;
wire  inst245_O;
wire  inst246_O;
wire  inst247_O;
wire  inst248_O;
wire  inst249_O;
wire  inst250_O;
wire  inst251_O;
wire  inst252_O;
wire  inst253_O;
wire  inst254_O;
wire  inst255_O;
Decode8 inst0 (.I(I), .O(inst0_O));
Decode8 inst1 (.I(I), .O(inst1_O));
Decode8 inst2 (.I(I), .O(inst2_O));
Decode8 inst3 (.I(I), .O(inst3_O));
Decode8 inst4 (.I(I), .O(inst4_O));
Decode8 inst5 (.I(I), .O(inst5_O));
Decode8 inst6 (.I(I), .O(inst6_O));
Decode8 inst7 (.I(I), .O(inst7_O));
Decode8 inst8 (.I(I), .O(inst8_O));
Decode8 inst9 (.I(I), .O(inst9_O));
Decode8 inst10 (.I(I), .O(inst10_O));
Decode8 inst11 (.I(I), .O(inst11_O));
Decode8 inst12 (.I(I), .O(inst12_O));
Decode8 inst13 (.I(I), .O(inst13_O));
Decode8 inst14 (.I(I), .O(inst14_O));
Decode8 inst15 (.I(I), .O(inst15_O));
Decode8 inst16 (.I(I), .O(inst16_O));
Decode8 inst17 (.I(I), .O(inst17_O));
Decode8 inst18 (.I(I), .O(inst18_O));
Decode8 inst19 (.I(I), .O(inst19_O));
Decode8 inst20 (.I(I), .O(inst20_O));
Decode8 inst21 (.I(I), .O(inst21_O));
Decode8 inst22 (.I(I), .O(inst22_O));
Decode8 inst23 (.I(I), .O(inst23_O));
Decode8 inst24 (.I(I), .O(inst24_O));
Decode8 inst25 (.I(I), .O(inst25_O));
Decode8 inst26 (.I(I), .O(inst26_O));
Decode8 inst27 (.I(I), .O(inst27_O));
Decode8 inst28 (.I(I), .O(inst28_O));
Decode8 inst29 (.I(I), .O(inst29_O));
Decode8 inst30 (.I(I), .O(inst30_O));
Decode8 inst31 (.I(I), .O(inst31_O));
Decode8 inst32 (.I(I), .O(inst32_O));
Decode8 inst33 (.I(I), .O(inst33_O));
Decode8 inst34 (.I(I), .O(inst34_O));
Decode8 inst35 (.I(I), .O(inst35_O));
Decode8 inst36 (.I(I), .O(inst36_O));
Decode8 inst37 (.I(I), .O(inst37_O));
Decode8 inst38 (.I(I), .O(inst38_O));
Decode8 inst39 (.I(I), .O(inst39_O));
Decode8 inst40 (.I(I), .O(inst40_O));
Decode8 inst41 (.I(I), .O(inst41_O));
Decode8 inst42 (.I(I), .O(inst42_O));
Decode8 inst43 (.I(I), .O(inst43_O));
Decode8 inst44 (.I(I), .O(inst44_O));
Decode8 inst45 (.I(I), .O(inst45_O));
Decode8 inst46 (.I(I), .O(inst46_O));
Decode8 inst47 (.I(I), .O(inst47_O));
Decode8 inst48 (.I(I), .O(inst48_O));
Decode8 inst49 (.I(I), .O(inst49_O));
Decode8 inst50 (.I(I), .O(inst50_O));
Decode8 inst51 (.I(I), .O(inst51_O));
Decode8 inst52 (.I(I), .O(inst52_O));
Decode8 inst53 (.I(I), .O(inst53_O));
Decode8 inst54 (.I(I), .O(inst54_O));
Decode8 inst55 (.I(I), .O(inst55_O));
Decode8 inst56 (.I(I), .O(inst56_O));
Decode8 inst57 (.I(I), .O(inst57_O));
Decode8 inst58 (.I(I), .O(inst58_O));
Decode8 inst59 (.I(I), .O(inst59_O));
Decode8 inst60 (.I(I), .O(inst60_O));
Decode8 inst61 (.I(I), .O(inst61_O));
Decode8 inst62 (.I(I), .O(inst62_O));
Decode8 inst63 (.I(I), .O(inst63_O));
Decode8 inst64 (.I(I), .O(inst64_O));
Decode8 inst65 (.I(I), .O(inst65_O));
Decode8 inst66 (.I(I), .O(inst66_O));
Decode8 inst67 (.I(I), .O(inst67_O));
Decode8 inst68 (.I(I), .O(inst68_O));
Decode8 inst69 (.I(I), .O(inst69_O));
Decode8 inst70 (.I(I), .O(inst70_O));
Decode8 inst71 (.I(I), .O(inst71_O));
Decode8 inst72 (.I(I), .O(inst72_O));
Decode8 inst73 (.I(I), .O(inst73_O));
Decode8 inst74 (.I(I), .O(inst74_O));
Decode8 inst75 (.I(I), .O(inst75_O));
Decode8 inst76 (.I(I), .O(inst76_O));
Decode8 inst77 (.I(I), .O(inst77_O));
Decode8 inst78 (.I(I), .O(inst78_O));
Decode8 inst79 (.I(I), .O(inst79_O));
Decode8 inst80 (.I(I), .O(inst80_O));
Decode8 inst81 (.I(I), .O(inst81_O));
Decode8 inst82 (.I(I), .O(inst82_O));
Decode8 inst83 (.I(I), .O(inst83_O));
Decode8 inst84 (.I(I), .O(inst84_O));
Decode8 inst85 (.I(I), .O(inst85_O));
Decode8 inst86 (.I(I), .O(inst86_O));
Decode8 inst87 (.I(I), .O(inst87_O));
Decode8 inst88 (.I(I), .O(inst88_O));
Decode8 inst89 (.I(I), .O(inst89_O));
Decode8 inst90 (.I(I), .O(inst90_O));
Decode8 inst91 (.I(I), .O(inst91_O));
Decode8 inst92 (.I(I), .O(inst92_O));
Decode8 inst93 (.I(I), .O(inst93_O));
Decode8 inst94 (.I(I), .O(inst94_O));
Decode8 inst95 (.I(I), .O(inst95_O));
Decode8 inst96 (.I(I), .O(inst96_O));
Decode8 inst97 (.I(I), .O(inst97_O));
Decode8 inst98 (.I(I), .O(inst98_O));
Decode8 inst99 (.I(I), .O(inst99_O));
Decode8 inst100 (.I(I), .O(inst100_O));
Decode8 inst101 (.I(I), .O(inst101_O));
Decode8 inst102 (.I(I), .O(inst102_O));
Decode8 inst103 (.I(I), .O(inst103_O));
Decode8 inst104 (.I(I), .O(inst104_O));
Decode8 inst105 (.I(I), .O(inst105_O));
Decode8 inst106 (.I(I), .O(inst106_O));
Decode8 inst107 (.I(I), .O(inst107_O));
Decode8 inst108 (.I(I), .O(inst108_O));
Decode8 inst109 (.I(I), .O(inst109_O));
Decode8 inst110 (.I(I), .O(inst110_O));
Decode8 inst111 (.I(I), .O(inst111_O));
Decode8 inst112 (.I(I), .O(inst112_O));
Decode8 inst113 (.I(I), .O(inst113_O));
Decode8 inst114 (.I(I), .O(inst114_O));
Decode8 inst115 (.I(I), .O(inst115_O));
Decode8 inst116 (.I(I), .O(inst116_O));
Decode8 inst117 (.I(I), .O(inst117_O));
Decode8 inst118 (.I(I), .O(inst118_O));
Decode8 inst119 (.I(I), .O(inst119_O));
Decode8 inst120 (.I(I), .O(inst120_O));
Decode8 inst121 (.I(I), .O(inst121_O));
Decode8 inst122 (.I(I), .O(inst122_O));
Decode8 inst123 (.I(I), .O(inst123_O));
Decode8 inst124 (.I(I), .O(inst124_O));
Decode8 inst125 (.I(I), .O(inst125_O));
Decode8 inst126 (.I(I), .O(inst126_O));
Decode8 inst127 (.I(I), .O(inst127_O));
Decode8 inst128 (.I(I), .O(inst128_O));
Decode8 inst129 (.I(I), .O(inst129_O));
Decode8 inst130 (.I(I), .O(inst130_O));
Decode8 inst131 (.I(I), .O(inst131_O));
Decode8 inst132 (.I(I), .O(inst132_O));
Decode8 inst133 (.I(I), .O(inst133_O));
Decode8 inst134 (.I(I), .O(inst134_O));
Decode8 inst135 (.I(I), .O(inst135_O));
Decode8 inst136 (.I(I), .O(inst136_O));
Decode8 inst137 (.I(I), .O(inst137_O));
Decode8 inst138 (.I(I), .O(inst138_O));
Decode8 inst139 (.I(I), .O(inst139_O));
Decode8 inst140 (.I(I), .O(inst140_O));
Decode8 inst141 (.I(I), .O(inst141_O));
Decode8 inst142 (.I(I), .O(inst142_O));
Decode8 inst143 (.I(I), .O(inst143_O));
Decode8 inst144 (.I(I), .O(inst144_O));
Decode8 inst145 (.I(I), .O(inst145_O));
Decode8 inst146 (.I(I), .O(inst146_O));
Decode8 inst147 (.I(I), .O(inst147_O));
Decode8 inst148 (.I(I), .O(inst148_O));
Decode8 inst149 (.I(I), .O(inst149_O));
Decode8 inst150 (.I(I), .O(inst150_O));
Decode8 inst151 (.I(I), .O(inst151_O));
Decode8 inst152 (.I(I), .O(inst152_O));
Decode8 inst153 (.I(I), .O(inst153_O));
Decode8 inst154 (.I(I), .O(inst154_O));
Decode8 inst155 (.I(I), .O(inst155_O));
Decode8 inst156 (.I(I), .O(inst156_O));
Decode8 inst157 (.I(I), .O(inst157_O));
Decode8 inst158 (.I(I), .O(inst158_O));
Decode8 inst159 (.I(I), .O(inst159_O));
Decode8 inst160 (.I(I), .O(inst160_O));
Decode8 inst161 (.I(I), .O(inst161_O));
Decode8 inst162 (.I(I), .O(inst162_O));
Decode8 inst163 (.I(I), .O(inst163_O));
Decode8 inst164 (.I(I), .O(inst164_O));
Decode8 inst165 (.I(I), .O(inst165_O));
Decode8 inst166 (.I(I), .O(inst166_O));
Decode8 inst167 (.I(I), .O(inst167_O));
Decode8 inst168 (.I(I), .O(inst168_O));
Decode8 inst169 (.I(I), .O(inst169_O));
Decode8 inst170 (.I(I), .O(inst170_O));
Decode8 inst171 (.I(I), .O(inst171_O));
Decode8 inst172 (.I(I), .O(inst172_O));
Decode8 inst173 (.I(I), .O(inst173_O));
Decode8 inst174 (.I(I), .O(inst174_O));
Decode8 inst175 (.I(I), .O(inst175_O));
Decode8 inst176 (.I(I), .O(inst176_O));
Decode8 inst177 (.I(I), .O(inst177_O));
Decode8 inst178 (.I(I), .O(inst178_O));
Decode8 inst179 (.I(I), .O(inst179_O));
Decode8 inst180 (.I(I), .O(inst180_O));
Decode8 inst181 (.I(I), .O(inst181_O));
Decode8 inst182 (.I(I), .O(inst182_O));
Decode8 inst183 (.I(I), .O(inst183_O));
Decode8 inst184 (.I(I), .O(inst184_O));
Decode8 inst185 (.I(I), .O(inst185_O));
Decode8 inst186 (.I(I), .O(inst186_O));
Decode8 inst187 (.I(I), .O(inst187_O));
Decode8 inst188 (.I(I), .O(inst188_O));
Decode8 inst189 (.I(I), .O(inst189_O));
Decode8 inst190 (.I(I), .O(inst190_O));
Decode8 inst191 (.I(I), .O(inst191_O));
Decode8 inst192 (.I(I), .O(inst192_O));
Decode8 inst193 (.I(I), .O(inst193_O));
Decode8 inst194 (.I(I), .O(inst194_O));
Decode8 inst195 (.I(I), .O(inst195_O));
Decode8 inst196 (.I(I), .O(inst196_O));
Decode8 inst197 (.I(I), .O(inst197_O));
Decode8 inst198 (.I(I), .O(inst198_O));
Decode8 inst199 (.I(I), .O(inst199_O));
Decode8 inst200 (.I(I), .O(inst200_O));
Decode8 inst201 (.I(I), .O(inst201_O));
Decode8 inst202 (.I(I), .O(inst202_O));
Decode8 inst203 (.I(I), .O(inst203_O));
Decode8 inst204 (.I(I), .O(inst204_O));
Decode8 inst205 (.I(I), .O(inst205_O));
Decode8 inst206 (.I(I), .O(inst206_O));
Decode8 inst207 (.I(I), .O(inst207_O));
Decode8 inst208 (.I(I), .O(inst208_O));
Decode8 inst209 (.I(I), .O(inst209_O));
Decode8 inst210 (.I(I), .O(inst210_O));
Decode8 inst211 (.I(I), .O(inst211_O));
Decode8 inst212 (.I(I), .O(inst212_O));
Decode8 inst213 (.I(I), .O(inst213_O));
Decode8 inst214 (.I(I), .O(inst214_O));
Decode8 inst215 (.I(I), .O(inst215_O));
Decode8 inst216 (.I(I), .O(inst216_O));
Decode8 inst217 (.I(I), .O(inst217_O));
Decode8 inst218 (.I(I), .O(inst218_O));
Decode8 inst219 (.I(I), .O(inst219_O));
Decode8 inst220 (.I(I), .O(inst220_O));
Decode8 inst221 (.I(I), .O(inst221_O));
Decode8 inst222 (.I(I), .O(inst222_O));
Decode8 inst223 (.I(I), .O(inst223_O));
Decode8 inst224 (.I(I), .O(inst224_O));
Decode8 inst225 (.I(I), .O(inst225_O));
Decode8 inst226 (.I(I), .O(inst226_O));
Decode8 inst227 (.I(I), .O(inst227_O));
Decode8 inst228 (.I(I), .O(inst228_O));
Decode8 inst229 (.I(I), .O(inst229_O));
Decode8 inst230 (.I(I), .O(inst230_O));
Decode8 inst231 (.I(I), .O(inst231_O));
Decode8 inst232 (.I(I), .O(inst232_O));
Decode8 inst233 (.I(I), .O(inst233_O));
Decode8 inst234 (.I(I), .O(inst234_O));
Decode8 inst235 (.I(I), .O(inst235_O));
Decode8 inst236 (.I(I), .O(inst236_O));
Decode8 inst237 (.I(I), .O(inst237_O));
Decode8 inst238 (.I(I), .O(inst238_O));
Decode8 inst239 (.I(I), .O(inst239_O));
Decode8 inst240 (.I(I), .O(inst240_O));
Decode8 inst241 (.I(I), .O(inst241_O));
Decode8 inst242 (.I(I), .O(inst242_O));
Decode8 inst243 (.I(I), .O(inst243_O));
Decode8 inst244 (.I(I), .O(inst244_O));
Decode8 inst245 (.I(I), .O(inst245_O));
Decode8 inst246 (.I(I), .O(inst246_O));
Decode8 inst247 (.I(I), .O(inst247_O));
Decode8 inst248 (.I(I), .O(inst248_O));
Decode8 inst249 (.I(I), .O(inst249_O));
Decode8 inst250 (.I(I), .O(inst250_O));
Decode8 inst251 (.I(I), .O(inst251_O));
Decode8 inst252 (.I(I), .O(inst252_O));
Decode8 inst253 (.I(I), .O(inst253_O));
Decode8 inst254 (.I(I), .O(inst254_O));
Decode8 inst255 (.I(I), .O(inst255_O));
assign O = {inst255_O,inst254_O,inst253_O,inst252_O,inst251_O,inst250_O,inst249_O,inst248_O,inst247_O,inst246_O,inst245_O,inst244_O,inst243_O,inst242_O,inst241_O,inst240_O,inst239_O,inst238_O,inst237_O,inst236_O,inst235_O,inst234_O,inst233_O,inst232_O,inst231_O,inst230_O,inst229_O,inst228_O,inst227_O,inst226_O,inst225_O,inst224_O,inst223_O,inst222_O,inst221_O,inst220_O,inst219_O,inst218_O,inst217_O,inst216_O,inst215_O,inst214_O,inst213_O,inst212_O,inst211_O,inst210_O,inst209_O,inst208_O,inst207_O,inst206_O,inst205_O,inst204_O,inst203_O,inst202_O,inst201_O,inst200_O,inst199_O,inst198_O,inst197_O,inst196_O,inst195_O,inst194_O,inst193_O,inst192_O,inst191_O,inst190_O,inst189_O,inst188_O,inst187_O,inst186_O,inst185_O,inst184_O,inst183_O,inst182_O,inst181_O,inst180_O,inst179_O,inst178_O,inst177_O,inst176_O,inst175_O,inst174_O,inst173_O,inst172_O,inst171_O,inst170_O,inst169_O,inst168_O,inst167_O,inst166_O,inst165_O,inst164_O,inst163_O,inst162_O,inst161_O,inst160_O,inst159_O,inst158_O,inst157_O,inst156_O,inst155_O,inst154_O,inst153_O,inst152_O,inst151_O,inst150_O,inst149_O,inst148_O,inst147_O,inst146_O,inst145_O,inst144_O,inst143_O,inst142_O,inst141_O,inst140_O,inst139_O,inst138_O,inst137_O,inst136_O,inst135_O,inst134_O,inst133_O,inst132_O,inst131_O,inst130_O,inst129_O,inst128_O,inst127_O,inst126_O,inst125_O,inst124_O,inst123_O,inst122_O,inst121_O,inst120_O,inst119_O,inst118_O,inst117_O,inst116_O,inst115_O,inst114_O,inst113_O,inst112_O,inst111_O,inst110_O,inst109_O,inst108_O,inst107_O,inst106_O,inst105_O,inst104_O,inst103_O,inst102_O,inst101_O,inst100_O,inst99_O,inst98_O,inst97_O,inst96_O,inst95_O,inst94_O,inst93_O,inst92_O,inst91_O,inst90_O,inst89_O,inst88_O,inst87_O,inst86_O,inst85_O,inst84_O,inst83_O,inst82_O,inst81_O,inst80_O,inst79_O,inst78_O,inst77_O,inst76_O,inst75_O,inst74_O,inst73_O,inst72_O,inst71_O,inst70_O,inst69_O,inst68_O,inst67_O,inst66_O,inst65_O,inst64_O,inst63_O,inst62_O,inst61_O,inst60_O,inst59_O,inst58_O,inst57_O,inst56_O,inst55_O,inst54_O,inst53_O,inst52_O,inst51_O,inst50_O,inst49_O,inst48_O,inst47_O,inst46_O,inst45_O,inst44_O,inst43_O,inst42_O,inst41_O,inst40_O,inst39_O,inst38_O,inst37_O,inst36_O,inst35_O,inst34_O,inst33_O,inst32_O,inst31_O,inst30_O,inst29_O,inst28_O,inst27_O,inst26_O,inst25_O,inst24_O,inst23_O,inst22_O,inst21_O,inst20_O,inst19_O,inst18_O,inst17_O,inst16_O,inst15_O,inst14_O,inst13_O,inst12_O,inst11_O,inst10_O,inst9_O,inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

