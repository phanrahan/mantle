module FixedLSR2_2 (input [1:0] I, output [1:0] O);
assign O = {1'b0,1'b0};
endmodule

