module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk, input [width-1:0] in, output [width-1:0] out);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module reg_P_wrapped (input CLK, input [7:0] I, output [7:0] O);
coreir_reg #(.clk_posedge(1'b1), .init(8'h00), .width(8)) reg_P_inst0(.clk(CLK), .in(I), .out(O));
endmodule

