module main (output  O, input  CLKIN);
wire  inst0_PLLOUTCORE;
wire  inst0_PLLOUTGLOBAL;
SB_PLL40_CORE #(.DIVF(7'b0111111),
.DIVQ(3'b101),
.DIVR(4'b0000),
.FEEDBACK_PATH("SIMPLE"),
.FILTER_RANGE(3'b001),
.PLLOUT_SELECT("GENCLK")) inst0 (.REFERENCECLK(CLKIN), .RESETB(1'b1), .BYPASS(1'b0), .PLLOUTCORE(inst0_PLLOUTCORE), .PLLOUTGLOBAL(inst0_PLLOUTGLOBAL));
assign O = inst0_PLLOUTGLOBAL;
endmodule

