module EQ8 (input [7:0] I0, input [7:0] I1, output  O);
wire  inst0_out;
coreir_eq inst0 (.in0(I0), .in1(I1), .out(inst0_out));
assign O = inst0_out;
endmodule

module Decode08 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode18 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode28 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode38 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode48 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode58 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode68 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode78 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode88 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode98 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode108 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode118 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode128 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode138 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode148 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode158 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode168 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode178 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode188 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode198 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode208 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode218 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode228 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode238 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode248 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode258 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode268 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode278 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode288 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode298 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode308 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode318 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode328 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode338 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode348 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode358 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode368 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode378 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode388 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode398 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode408 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode418 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode428 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode438 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode448 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode458 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode468 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode478 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode488 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode498 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode508 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode518 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode528 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode538 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode548 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode558 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode568 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode578 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode588 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode598 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode608 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode618 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode628 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode638 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode648 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode658 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode668 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode678 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode688 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode698 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode708 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode718 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode728 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode738 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode748 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode758 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode768 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode778 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode788 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode798 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode808 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode818 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode828 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode838 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode848 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode858 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode868 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode878 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode888 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode898 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode908 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode918 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode928 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode938 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode948 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode958 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode968 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode978 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode988 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode998 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1008 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1018 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1028 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1038 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1048 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1058 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1068 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1078 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1088 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1098 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1108 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1118 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1128 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1138 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1148 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1158 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1168 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1178 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1188 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1198 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1208 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1218 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1228 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1238 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1248 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1258 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1268 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1278 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1288 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1298 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1308 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1318 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1328 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1338 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1348 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1358 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1368 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1378 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1388 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1398 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1408 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1418 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1428 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1438 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1448 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1458 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1468 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1478 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1488 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1498 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1508 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1518 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1528 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1538 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1548 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1558 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1568 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1578 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1588 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1598 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1608 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1618 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1628 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1638 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1648 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1658 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1668 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1678 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1688 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1698 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1708 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1718 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1728 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1738 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1748 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1758 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1768 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1778 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1788 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1798 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1808 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1818 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1828 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1838 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1848 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1858 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1868 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1878 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1888 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1898 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1908 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1918 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1928 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1938 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1948 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1958 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1968 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1978 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1988 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode1998 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2008 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2018 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2028 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2038 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2048 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2058 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2068 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2078 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2088 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2098 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2108 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2118 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2128 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2138 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2148 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2158 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2168 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2178 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2188 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2198 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2208 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2218 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2228 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2238 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2248 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2258 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2268 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2278 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2288 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2298 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2308 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2318 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2328 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2338 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2348 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2358 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2368 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2378 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2388 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2398 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2408 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2418 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2428 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2438 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2448 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2458 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2468 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2478 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2488 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2498 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2508 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2518 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2528 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2538 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2548 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decode2558 (input [7:0] I, output  O);
wire  inst0_O;
EQ8 inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
assign O = inst0_O;
endmodule

module Decoder8 (input [7:0] I, output [255:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
wire  inst64_O;
wire  inst65_O;
wire  inst66_O;
wire  inst67_O;
wire  inst68_O;
wire  inst69_O;
wire  inst70_O;
wire  inst71_O;
wire  inst72_O;
wire  inst73_O;
wire  inst74_O;
wire  inst75_O;
wire  inst76_O;
wire  inst77_O;
wire  inst78_O;
wire  inst79_O;
wire  inst80_O;
wire  inst81_O;
wire  inst82_O;
wire  inst83_O;
wire  inst84_O;
wire  inst85_O;
wire  inst86_O;
wire  inst87_O;
wire  inst88_O;
wire  inst89_O;
wire  inst90_O;
wire  inst91_O;
wire  inst92_O;
wire  inst93_O;
wire  inst94_O;
wire  inst95_O;
wire  inst96_O;
wire  inst97_O;
wire  inst98_O;
wire  inst99_O;
wire  inst100_O;
wire  inst101_O;
wire  inst102_O;
wire  inst103_O;
wire  inst104_O;
wire  inst105_O;
wire  inst106_O;
wire  inst107_O;
wire  inst108_O;
wire  inst109_O;
wire  inst110_O;
wire  inst111_O;
wire  inst112_O;
wire  inst113_O;
wire  inst114_O;
wire  inst115_O;
wire  inst116_O;
wire  inst117_O;
wire  inst118_O;
wire  inst119_O;
wire  inst120_O;
wire  inst121_O;
wire  inst122_O;
wire  inst123_O;
wire  inst124_O;
wire  inst125_O;
wire  inst126_O;
wire  inst127_O;
wire  inst128_O;
wire  inst129_O;
wire  inst130_O;
wire  inst131_O;
wire  inst132_O;
wire  inst133_O;
wire  inst134_O;
wire  inst135_O;
wire  inst136_O;
wire  inst137_O;
wire  inst138_O;
wire  inst139_O;
wire  inst140_O;
wire  inst141_O;
wire  inst142_O;
wire  inst143_O;
wire  inst144_O;
wire  inst145_O;
wire  inst146_O;
wire  inst147_O;
wire  inst148_O;
wire  inst149_O;
wire  inst150_O;
wire  inst151_O;
wire  inst152_O;
wire  inst153_O;
wire  inst154_O;
wire  inst155_O;
wire  inst156_O;
wire  inst157_O;
wire  inst158_O;
wire  inst159_O;
wire  inst160_O;
wire  inst161_O;
wire  inst162_O;
wire  inst163_O;
wire  inst164_O;
wire  inst165_O;
wire  inst166_O;
wire  inst167_O;
wire  inst168_O;
wire  inst169_O;
wire  inst170_O;
wire  inst171_O;
wire  inst172_O;
wire  inst173_O;
wire  inst174_O;
wire  inst175_O;
wire  inst176_O;
wire  inst177_O;
wire  inst178_O;
wire  inst179_O;
wire  inst180_O;
wire  inst181_O;
wire  inst182_O;
wire  inst183_O;
wire  inst184_O;
wire  inst185_O;
wire  inst186_O;
wire  inst187_O;
wire  inst188_O;
wire  inst189_O;
wire  inst190_O;
wire  inst191_O;
wire  inst192_O;
wire  inst193_O;
wire  inst194_O;
wire  inst195_O;
wire  inst196_O;
wire  inst197_O;
wire  inst198_O;
wire  inst199_O;
wire  inst200_O;
wire  inst201_O;
wire  inst202_O;
wire  inst203_O;
wire  inst204_O;
wire  inst205_O;
wire  inst206_O;
wire  inst207_O;
wire  inst208_O;
wire  inst209_O;
wire  inst210_O;
wire  inst211_O;
wire  inst212_O;
wire  inst213_O;
wire  inst214_O;
wire  inst215_O;
wire  inst216_O;
wire  inst217_O;
wire  inst218_O;
wire  inst219_O;
wire  inst220_O;
wire  inst221_O;
wire  inst222_O;
wire  inst223_O;
wire  inst224_O;
wire  inst225_O;
wire  inst226_O;
wire  inst227_O;
wire  inst228_O;
wire  inst229_O;
wire  inst230_O;
wire  inst231_O;
wire  inst232_O;
wire  inst233_O;
wire  inst234_O;
wire  inst235_O;
wire  inst236_O;
wire  inst237_O;
wire  inst238_O;
wire  inst239_O;
wire  inst240_O;
wire  inst241_O;
wire  inst242_O;
wire  inst243_O;
wire  inst244_O;
wire  inst245_O;
wire  inst246_O;
wire  inst247_O;
wire  inst248_O;
wire  inst249_O;
wire  inst250_O;
wire  inst251_O;
wire  inst252_O;
wire  inst253_O;
wire  inst254_O;
wire  inst255_O;
Decode08 inst0 (.I(I), .O(inst0_O));
Decode18 inst1 (.I(I), .O(inst1_O));
Decode28 inst2 (.I(I), .O(inst2_O));
Decode38 inst3 (.I(I), .O(inst3_O));
Decode48 inst4 (.I(I), .O(inst4_O));
Decode58 inst5 (.I(I), .O(inst5_O));
Decode68 inst6 (.I(I), .O(inst6_O));
Decode78 inst7 (.I(I), .O(inst7_O));
Decode88 inst8 (.I(I), .O(inst8_O));
Decode98 inst9 (.I(I), .O(inst9_O));
Decode108 inst10 (.I(I), .O(inst10_O));
Decode118 inst11 (.I(I), .O(inst11_O));
Decode128 inst12 (.I(I), .O(inst12_O));
Decode138 inst13 (.I(I), .O(inst13_O));
Decode148 inst14 (.I(I), .O(inst14_O));
Decode158 inst15 (.I(I), .O(inst15_O));
Decode168 inst16 (.I(I), .O(inst16_O));
Decode178 inst17 (.I(I), .O(inst17_O));
Decode188 inst18 (.I(I), .O(inst18_O));
Decode198 inst19 (.I(I), .O(inst19_O));
Decode208 inst20 (.I(I), .O(inst20_O));
Decode218 inst21 (.I(I), .O(inst21_O));
Decode228 inst22 (.I(I), .O(inst22_O));
Decode238 inst23 (.I(I), .O(inst23_O));
Decode248 inst24 (.I(I), .O(inst24_O));
Decode258 inst25 (.I(I), .O(inst25_O));
Decode268 inst26 (.I(I), .O(inst26_O));
Decode278 inst27 (.I(I), .O(inst27_O));
Decode288 inst28 (.I(I), .O(inst28_O));
Decode298 inst29 (.I(I), .O(inst29_O));
Decode308 inst30 (.I(I), .O(inst30_O));
Decode318 inst31 (.I(I), .O(inst31_O));
Decode328 inst32 (.I(I), .O(inst32_O));
Decode338 inst33 (.I(I), .O(inst33_O));
Decode348 inst34 (.I(I), .O(inst34_O));
Decode358 inst35 (.I(I), .O(inst35_O));
Decode368 inst36 (.I(I), .O(inst36_O));
Decode378 inst37 (.I(I), .O(inst37_O));
Decode388 inst38 (.I(I), .O(inst38_O));
Decode398 inst39 (.I(I), .O(inst39_O));
Decode408 inst40 (.I(I), .O(inst40_O));
Decode418 inst41 (.I(I), .O(inst41_O));
Decode428 inst42 (.I(I), .O(inst42_O));
Decode438 inst43 (.I(I), .O(inst43_O));
Decode448 inst44 (.I(I), .O(inst44_O));
Decode458 inst45 (.I(I), .O(inst45_O));
Decode468 inst46 (.I(I), .O(inst46_O));
Decode478 inst47 (.I(I), .O(inst47_O));
Decode488 inst48 (.I(I), .O(inst48_O));
Decode498 inst49 (.I(I), .O(inst49_O));
Decode508 inst50 (.I(I), .O(inst50_O));
Decode518 inst51 (.I(I), .O(inst51_O));
Decode528 inst52 (.I(I), .O(inst52_O));
Decode538 inst53 (.I(I), .O(inst53_O));
Decode548 inst54 (.I(I), .O(inst54_O));
Decode558 inst55 (.I(I), .O(inst55_O));
Decode568 inst56 (.I(I), .O(inst56_O));
Decode578 inst57 (.I(I), .O(inst57_O));
Decode588 inst58 (.I(I), .O(inst58_O));
Decode598 inst59 (.I(I), .O(inst59_O));
Decode608 inst60 (.I(I), .O(inst60_O));
Decode618 inst61 (.I(I), .O(inst61_O));
Decode628 inst62 (.I(I), .O(inst62_O));
Decode638 inst63 (.I(I), .O(inst63_O));
Decode648 inst64 (.I(I), .O(inst64_O));
Decode658 inst65 (.I(I), .O(inst65_O));
Decode668 inst66 (.I(I), .O(inst66_O));
Decode678 inst67 (.I(I), .O(inst67_O));
Decode688 inst68 (.I(I), .O(inst68_O));
Decode698 inst69 (.I(I), .O(inst69_O));
Decode708 inst70 (.I(I), .O(inst70_O));
Decode718 inst71 (.I(I), .O(inst71_O));
Decode728 inst72 (.I(I), .O(inst72_O));
Decode738 inst73 (.I(I), .O(inst73_O));
Decode748 inst74 (.I(I), .O(inst74_O));
Decode758 inst75 (.I(I), .O(inst75_O));
Decode768 inst76 (.I(I), .O(inst76_O));
Decode778 inst77 (.I(I), .O(inst77_O));
Decode788 inst78 (.I(I), .O(inst78_O));
Decode798 inst79 (.I(I), .O(inst79_O));
Decode808 inst80 (.I(I), .O(inst80_O));
Decode818 inst81 (.I(I), .O(inst81_O));
Decode828 inst82 (.I(I), .O(inst82_O));
Decode838 inst83 (.I(I), .O(inst83_O));
Decode848 inst84 (.I(I), .O(inst84_O));
Decode858 inst85 (.I(I), .O(inst85_O));
Decode868 inst86 (.I(I), .O(inst86_O));
Decode878 inst87 (.I(I), .O(inst87_O));
Decode888 inst88 (.I(I), .O(inst88_O));
Decode898 inst89 (.I(I), .O(inst89_O));
Decode908 inst90 (.I(I), .O(inst90_O));
Decode918 inst91 (.I(I), .O(inst91_O));
Decode928 inst92 (.I(I), .O(inst92_O));
Decode938 inst93 (.I(I), .O(inst93_O));
Decode948 inst94 (.I(I), .O(inst94_O));
Decode958 inst95 (.I(I), .O(inst95_O));
Decode968 inst96 (.I(I), .O(inst96_O));
Decode978 inst97 (.I(I), .O(inst97_O));
Decode988 inst98 (.I(I), .O(inst98_O));
Decode998 inst99 (.I(I), .O(inst99_O));
Decode1008 inst100 (.I(I), .O(inst100_O));
Decode1018 inst101 (.I(I), .O(inst101_O));
Decode1028 inst102 (.I(I), .O(inst102_O));
Decode1038 inst103 (.I(I), .O(inst103_O));
Decode1048 inst104 (.I(I), .O(inst104_O));
Decode1058 inst105 (.I(I), .O(inst105_O));
Decode1068 inst106 (.I(I), .O(inst106_O));
Decode1078 inst107 (.I(I), .O(inst107_O));
Decode1088 inst108 (.I(I), .O(inst108_O));
Decode1098 inst109 (.I(I), .O(inst109_O));
Decode1108 inst110 (.I(I), .O(inst110_O));
Decode1118 inst111 (.I(I), .O(inst111_O));
Decode1128 inst112 (.I(I), .O(inst112_O));
Decode1138 inst113 (.I(I), .O(inst113_O));
Decode1148 inst114 (.I(I), .O(inst114_O));
Decode1158 inst115 (.I(I), .O(inst115_O));
Decode1168 inst116 (.I(I), .O(inst116_O));
Decode1178 inst117 (.I(I), .O(inst117_O));
Decode1188 inst118 (.I(I), .O(inst118_O));
Decode1198 inst119 (.I(I), .O(inst119_O));
Decode1208 inst120 (.I(I), .O(inst120_O));
Decode1218 inst121 (.I(I), .O(inst121_O));
Decode1228 inst122 (.I(I), .O(inst122_O));
Decode1238 inst123 (.I(I), .O(inst123_O));
Decode1248 inst124 (.I(I), .O(inst124_O));
Decode1258 inst125 (.I(I), .O(inst125_O));
Decode1268 inst126 (.I(I), .O(inst126_O));
Decode1278 inst127 (.I(I), .O(inst127_O));
Decode1288 inst128 (.I(I), .O(inst128_O));
Decode1298 inst129 (.I(I), .O(inst129_O));
Decode1308 inst130 (.I(I), .O(inst130_O));
Decode1318 inst131 (.I(I), .O(inst131_O));
Decode1328 inst132 (.I(I), .O(inst132_O));
Decode1338 inst133 (.I(I), .O(inst133_O));
Decode1348 inst134 (.I(I), .O(inst134_O));
Decode1358 inst135 (.I(I), .O(inst135_O));
Decode1368 inst136 (.I(I), .O(inst136_O));
Decode1378 inst137 (.I(I), .O(inst137_O));
Decode1388 inst138 (.I(I), .O(inst138_O));
Decode1398 inst139 (.I(I), .O(inst139_O));
Decode1408 inst140 (.I(I), .O(inst140_O));
Decode1418 inst141 (.I(I), .O(inst141_O));
Decode1428 inst142 (.I(I), .O(inst142_O));
Decode1438 inst143 (.I(I), .O(inst143_O));
Decode1448 inst144 (.I(I), .O(inst144_O));
Decode1458 inst145 (.I(I), .O(inst145_O));
Decode1468 inst146 (.I(I), .O(inst146_O));
Decode1478 inst147 (.I(I), .O(inst147_O));
Decode1488 inst148 (.I(I), .O(inst148_O));
Decode1498 inst149 (.I(I), .O(inst149_O));
Decode1508 inst150 (.I(I), .O(inst150_O));
Decode1518 inst151 (.I(I), .O(inst151_O));
Decode1528 inst152 (.I(I), .O(inst152_O));
Decode1538 inst153 (.I(I), .O(inst153_O));
Decode1548 inst154 (.I(I), .O(inst154_O));
Decode1558 inst155 (.I(I), .O(inst155_O));
Decode1568 inst156 (.I(I), .O(inst156_O));
Decode1578 inst157 (.I(I), .O(inst157_O));
Decode1588 inst158 (.I(I), .O(inst158_O));
Decode1598 inst159 (.I(I), .O(inst159_O));
Decode1608 inst160 (.I(I), .O(inst160_O));
Decode1618 inst161 (.I(I), .O(inst161_O));
Decode1628 inst162 (.I(I), .O(inst162_O));
Decode1638 inst163 (.I(I), .O(inst163_O));
Decode1648 inst164 (.I(I), .O(inst164_O));
Decode1658 inst165 (.I(I), .O(inst165_O));
Decode1668 inst166 (.I(I), .O(inst166_O));
Decode1678 inst167 (.I(I), .O(inst167_O));
Decode1688 inst168 (.I(I), .O(inst168_O));
Decode1698 inst169 (.I(I), .O(inst169_O));
Decode1708 inst170 (.I(I), .O(inst170_O));
Decode1718 inst171 (.I(I), .O(inst171_O));
Decode1728 inst172 (.I(I), .O(inst172_O));
Decode1738 inst173 (.I(I), .O(inst173_O));
Decode1748 inst174 (.I(I), .O(inst174_O));
Decode1758 inst175 (.I(I), .O(inst175_O));
Decode1768 inst176 (.I(I), .O(inst176_O));
Decode1778 inst177 (.I(I), .O(inst177_O));
Decode1788 inst178 (.I(I), .O(inst178_O));
Decode1798 inst179 (.I(I), .O(inst179_O));
Decode1808 inst180 (.I(I), .O(inst180_O));
Decode1818 inst181 (.I(I), .O(inst181_O));
Decode1828 inst182 (.I(I), .O(inst182_O));
Decode1838 inst183 (.I(I), .O(inst183_O));
Decode1848 inst184 (.I(I), .O(inst184_O));
Decode1858 inst185 (.I(I), .O(inst185_O));
Decode1868 inst186 (.I(I), .O(inst186_O));
Decode1878 inst187 (.I(I), .O(inst187_O));
Decode1888 inst188 (.I(I), .O(inst188_O));
Decode1898 inst189 (.I(I), .O(inst189_O));
Decode1908 inst190 (.I(I), .O(inst190_O));
Decode1918 inst191 (.I(I), .O(inst191_O));
Decode1928 inst192 (.I(I), .O(inst192_O));
Decode1938 inst193 (.I(I), .O(inst193_O));
Decode1948 inst194 (.I(I), .O(inst194_O));
Decode1958 inst195 (.I(I), .O(inst195_O));
Decode1968 inst196 (.I(I), .O(inst196_O));
Decode1978 inst197 (.I(I), .O(inst197_O));
Decode1988 inst198 (.I(I), .O(inst198_O));
Decode1998 inst199 (.I(I), .O(inst199_O));
Decode2008 inst200 (.I(I), .O(inst200_O));
Decode2018 inst201 (.I(I), .O(inst201_O));
Decode2028 inst202 (.I(I), .O(inst202_O));
Decode2038 inst203 (.I(I), .O(inst203_O));
Decode2048 inst204 (.I(I), .O(inst204_O));
Decode2058 inst205 (.I(I), .O(inst205_O));
Decode2068 inst206 (.I(I), .O(inst206_O));
Decode2078 inst207 (.I(I), .O(inst207_O));
Decode2088 inst208 (.I(I), .O(inst208_O));
Decode2098 inst209 (.I(I), .O(inst209_O));
Decode2108 inst210 (.I(I), .O(inst210_O));
Decode2118 inst211 (.I(I), .O(inst211_O));
Decode2128 inst212 (.I(I), .O(inst212_O));
Decode2138 inst213 (.I(I), .O(inst213_O));
Decode2148 inst214 (.I(I), .O(inst214_O));
Decode2158 inst215 (.I(I), .O(inst215_O));
Decode2168 inst216 (.I(I), .O(inst216_O));
Decode2178 inst217 (.I(I), .O(inst217_O));
Decode2188 inst218 (.I(I), .O(inst218_O));
Decode2198 inst219 (.I(I), .O(inst219_O));
Decode2208 inst220 (.I(I), .O(inst220_O));
Decode2218 inst221 (.I(I), .O(inst221_O));
Decode2228 inst222 (.I(I), .O(inst222_O));
Decode2238 inst223 (.I(I), .O(inst223_O));
Decode2248 inst224 (.I(I), .O(inst224_O));
Decode2258 inst225 (.I(I), .O(inst225_O));
Decode2268 inst226 (.I(I), .O(inst226_O));
Decode2278 inst227 (.I(I), .O(inst227_O));
Decode2288 inst228 (.I(I), .O(inst228_O));
Decode2298 inst229 (.I(I), .O(inst229_O));
Decode2308 inst230 (.I(I), .O(inst230_O));
Decode2318 inst231 (.I(I), .O(inst231_O));
Decode2328 inst232 (.I(I), .O(inst232_O));
Decode2338 inst233 (.I(I), .O(inst233_O));
Decode2348 inst234 (.I(I), .O(inst234_O));
Decode2358 inst235 (.I(I), .O(inst235_O));
Decode2368 inst236 (.I(I), .O(inst236_O));
Decode2378 inst237 (.I(I), .O(inst237_O));
Decode2388 inst238 (.I(I), .O(inst238_O));
Decode2398 inst239 (.I(I), .O(inst239_O));
Decode2408 inst240 (.I(I), .O(inst240_O));
Decode2418 inst241 (.I(I), .O(inst241_O));
Decode2428 inst242 (.I(I), .O(inst242_O));
Decode2438 inst243 (.I(I), .O(inst243_O));
Decode2448 inst244 (.I(I), .O(inst244_O));
Decode2458 inst245 (.I(I), .O(inst245_O));
Decode2468 inst246 (.I(I), .O(inst246_O));
Decode2478 inst247 (.I(I), .O(inst247_O));
Decode2488 inst248 (.I(I), .O(inst248_O));
Decode2498 inst249 (.I(I), .O(inst249_O));
Decode2508 inst250 (.I(I), .O(inst250_O));
Decode2518 inst251 (.I(I), .O(inst251_O));
Decode2528 inst252 (.I(I), .O(inst252_O));
Decode2538 inst253 (.I(I), .O(inst253_O));
Decode2548 inst254 (.I(I), .O(inst254_O));
Decode2558 inst255 (.I(I), .O(inst255_O));
assign O = {inst255_O,inst254_O,inst253_O,inst252_O,inst251_O,inst250_O,inst249_O,inst248_O,inst247_O,inst246_O,inst245_O,inst244_O,inst243_O,inst242_O,inst241_O,inst240_O,inst239_O,inst238_O,inst237_O,inst236_O,inst235_O,inst234_O,inst233_O,inst232_O,inst231_O,inst230_O,inst229_O,inst228_O,inst227_O,inst226_O,inst225_O,inst224_O,inst223_O,inst222_O,inst221_O,inst220_O,inst219_O,inst218_O,inst217_O,inst216_O,inst215_O,inst214_O,inst213_O,inst212_O,inst211_O,inst210_O,inst209_O,inst208_O,inst207_O,inst206_O,inst205_O,inst204_O,inst203_O,inst202_O,inst201_O,inst200_O,inst199_O,inst198_O,inst197_O,inst196_O,inst195_O,inst194_O,inst193_O,inst192_O,inst191_O,inst190_O,inst189_O,inst188_O,inst187_O,inst186_O,inst185_O,inst184_O,inst183_O,inst182_O,inst181_O,inst180_O,inst179_O,inst178_O,inst177_O,inst176_O,inst175_O,inst174_O,inst173_O,inst172_O,inst171_O,inst170_O,inst169_O,inst168_O,inst167_O,inst166_O,inst165_O,inst164_O,inst163_O,inst162_O,inst161_O,inst160_O,inst159_O,inst158_O,inst157_O,inst156_O,inst155_O,inst154_O,inst153_O,inst152_O,inst151_O,inst150_O,inst149_O,inst148_O,inst147_O,inst146_O,inst145_O,inst144_O,inst143_O,inst142_O,inst141_O,inst140_O,inst139_O,inst138_O,inst137_O,inst136_O,inst135_O,inst134_O,inst133_O,inst132_O,inst131_O,inst130_O,inst129_O,inst128_O,inst127_O,inst126_O,inst125_O,inst124_O,inst123_O,inst122_O,inst121_O,inst120_O,inst119_O,inst118_O,inst117_O,inst116_O,inst115_O,inst114_O,inst113_O,inst112_O,inst111_O,inst110_O,inst109_O,inst108_O,inst107_O,inst106_O,inst105_O,inst104_O,inst103_O,inst102_O,inst101_O,inst100_O,inst99_O,inst98_O,inst97_O,inst96_O,inst95_O,inst94_O,inst93_O,inst92_O,inst91_O,inst90_O,inst89_O,inst88_O,inst87_O,inst86_O,inst85_O,inst84_O,inst83_O,inst82_O,inst81_O,inst80_O,inst79_O,inst78_O,inst77_O,inst76_O,inst75_O,inst74_O,inst73_O,inst72_O,inst71_O,inst70_O,inst69_O,inst68_O,inst67_O,inst66_O,inst65_O,inst64_O,inst63_O,inst62_O,inst61_O,inst60_O,inst59_O,inst58_O,inst57_O,inst56_O,inst55_O,inst54_O,inst53_O,inst52_O,inst51_O,inst50_O,inst49_O,inst48_O,inst47_O,inst46_O,inst45_O,inst44_O,inst43_O,inst42_O,inst41_O,inst40_O,inst39_O,inst38_O,inst37_O,inst36_O,inst35_O,inst34_O,inst33_O,inst32_O,inst31_O,inst30_O,inst29_O,inst28_O,inst27_O,inst26_O,inst25_O,inst24_O,inst23_O,inst22_O,inst21_O,inst20_O,inst19_O,inst18_O,inst17_O,inst16_O,inst15_O,inst14_O,inst13_O,inst12_O,inst11_O,inst10_O,inst9_O,inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

