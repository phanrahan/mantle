module main (output [7:0] LED, input [7:0] SWITCH, input  CLKIN);
wire  inst0_DOA;
wire  inst0_DOB;
wire  inst0_DOC;
wire  inst0_DOD;
RAM64M #(.INIT_A(64'hAAAAAAAAAAAAAAAA),
.INIT_C(64'h5555555555555555),
.INIT_B(64'hFFFFFFFFFFFFFFFF),
.INIT_D(64'h0000000000000000)) inst0 (.ADDRA({SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .ADDRB({SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .ADDRC({SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .ADDRD({SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .DIA(1'b0), .DIB(1'b0), .DIC(1'b0), .DID(1'b0), .DOA(inst0_DOA), .DOB(inst0_DOB), .DOC(inst0_DOC), .DOD(inst0_DOD), .WE(1'b0), .WCLK(CLKIN));
assign LED = {inst0_DOD,inst0_DOD,inst0_DOC,inst0_DOC,inst0_DOB,inst0_DOB,inst0_DOA,inst0_DOA};
endmodule

