module main (input  I0, input  I1, input  I2, input  I3, input  I4, input  I5, input  I6, input  I7, output  D7, output  D6, output  D5, output  D4, output  D3, output  D2, output  D1, output  D0, input  CLKIN);
wire [15:0] inst0_RDATA;
SB_RAM40_4K #(.INIT_0(256'h000F000E000D000C000B000A0009000800070006000500040003000200010000),
.INIT_1(256'h001F001E001D001C001B001A0019001800170016001500140013001200110010),
.INIT_2(256'h002F002E002D002C002B002A0029002800270026002500240023002200210020),
.INIT_3(256'h003F003E003D003C003B003A0039003800370036003500340033003200310030),
.INIT_4(256'h004F004E004D004C004B004A0049004800470046004500440043004200410040),
.INIT_5(256'h005F005E005D005C005B005A0059005800570056005500540053005200510050),
.INIT_6(256'h006F006E006D006C006B006A0069006800670066006500640063006200610060),
.INIT_7(256'h007F007E007D007C007B007A0079007800770076007500740073007200710070),
.INIT_8(256'h008F008E008D008C008B008A0089008800870086008500840083008200810080),
.INIT_9(256'h009F009E009D009C009B009A0099009800970096009500940093009200910090),
.INIT_A(256'h00AF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A0),
.INIT_B(256'h00BF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B0),
.INIT_C(256'h00CF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C0),
.INIT_D(256'h00DF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D0),
.INIT_E(256'h00EF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E0),
.INIT_F(256'h00FF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F0),
.READ_MODE(0),
.WRITE_MODE(0)) inst0 (.RDATA(inst0_RDATA), .RADDR({1'b0,1'b0,1'b0,I7,I6,I5,I4,I3,I2,I1,I0}), .RCLK(CLKIN), .RCLKE(1'b1), .RE(1'b1), .WCLK(CLKIN), .WCLKE(1'b0), .WE(1'b0), .WADDR({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .MASK({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .WDATA({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
assign D7 = inst0_RDATA[7];
assign D6 = inst0_RDATA[6];
assign D5 = inst0_RDATA[5];
assign D4 = inst0_RDATA[4];
assign D3 = inst0_RDATA[3];
assign D2 = inst0_RDATA[2];
assign D1 = inst0_RDATA[1];
assign D0 = inst0_RDATA[0];
endmodule

