module FixedLSL4_0 (input [3:0] I, output [3:0] O);
assign O = I;
endmodule

