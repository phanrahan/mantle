module Adders8_6_8_cinNone_coutNone (input [7:0] I0, input [7:0] I1, output [7:0] O);
wire  inst0_O;
wire  inst1_LO;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_LO;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_LO;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_LO;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_LO;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_LO;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_LO;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_LO;
wire  inst30_O;
wire  inst31_O;
LUT2 #(.INIT(4'h6)) inst0 (.I0(I0[0]), .I1(I1[0]), .O(inst0_O));
MULT_AND inst1 (.I0(I0[0]), .I1(I1[0]), .LO(inst1_LO));
MUXCY inst2 (.DI(inst1_LO), .CI(1'b0), .S(inst0_O), .O(inst2_O));
XORCY inst3 (.LI(inst0_O), .CI(1'b0), .O(inst3_O));
LUT2 #(.INIT(4'h6)) inst4 (.I0(I0[1]), .I1(I1[1]), .O(inst4_O));
MULT_AND inst5 (.I0(I0[1]), .I1(I1[1]), .LO(inst5_LO));
MUXCY inst6 (.DI(inst5_LO), .CI(inst2_O), .S(inst4_O), .O(inst6_O));
XORCY inst7 (.LI(inst4_O), .CI(inst2_O), .O(inst7_O));
LUT2 #(.INIT(4'h6)) inst8 (.I0(I0[2]), .I1(I1[2]), .O(inst8_O));
MULT_AND inst9 (.I0(I0[2]), .I1(I1[2]), .LO(inst9_LO));
MUXCY inst10 (.DI(inst9_LO), .CI(inst6_O), .S(inst8_O), .O(inst10_O));
XORCY inst11 (.LI(inst8_O), .CI(inst6_O), .O(inst11_O));
LUT2 #(.INIT(4'h6)) inst12 (.I0(I0[3]), .I1(I1[3]), .O(inst12_O));
MULT_AND inst13 (.I0(I0[3]), .I1(I1[3]), .LO(inst13_LO));
MUXCY inst14 (.DI(inst13_LO), .CI(inst10_O), .S(inst12_O), .O(inst14_O));
XORCY inst15 (.LI(inst12_O), .CI(inst10_O), .O(inst15_O));
LUT2 #(.INIT(4'h6)) inst16 (.I0(I0[4]), .I1(I1[4]), .O(inst16_O));
MULT_AND inst17 (.I0(I0[4]), .I1(I1[4]), .LO(inst17_LO));
MUXCY inst18 (.DI(inst17_LO), .CI(inst14_O), .S(inst16_O), .O(inst18_O));
XORCY inst19 (.LI(inst16_O), .CI(inst14_O), .O(inst19_O));
LUT2 #(.INIT(4'h6)) inst20 (.I0(I0[5]), .I1(I1[5]), .O(inst20_O));
MULT_AND inst21 (.I0(I0[5]), .I1(I1[5]), .LO(inst21_LO));
MUXCY inst22 (.DI(inst21_LO), .CI(inst18_O), .S(inst20_O), .O(inst22_O));
XORCY inst23 (.LI(inst20_O), .CI(inst18_O), .O(inst23_O));
LUT2 #(.INIT(4'h6)) inst24 (.I0(I0[6]), .I1(I1[6]), .O(inst24_O));
MULT_AND inst25 (.I0(I0[6]), .I1(I1[6]), .LO(inst25_LO));
MUXCY inst26 (.DI(inst25_LO), .CI(inst22_O), .S(inst24_O), .O(inst26_O));
XORCY inst27 (.LI(inst24_O), .CI(inst22_O), .O(inst27_O));
LUT2 #(.INIT(4'h6)) inst28 (.I0(I0[7]), .I1(I1[7]), .O(inst28_O));
MULT_AND inst29 (.I0(I0[7]), .I1(I1[7]), .LO(inst29_LO));
MUXCY inst30 (.DI(inst29_LO), .CI(inst26_O), .S(inst28_O), .O(inst30_O));
XORCY inst31 (.LI(inst28_O), .CI(inst26_O), .O(inst31_O));
assign O = {inst31_O,inst27_O,inst23_O,inst19_O,inst15_O,inst11_O,inst7_O,inst3_O};
endmodule

module Arbiter8 (input [7:0] I, output [7:0] O);
wire [7:0] inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
Adders8_6_8_cinNone_coutNone inst0 (.I0(I), .I1({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst0_O));
LUT2 #(.INIT(4'h2)) inst1 (.I0(I[0]), .I1(inst0_O[0]), .O(inst1_O));
LUT2 #(.INIT(4'h2)) inst2 (.I0(I[1]), .I1(inst0_O[1]), .O(inst2_O));
LUT2 #(.INIT(4'h2)) inst3 (.I0(I[2]), .I1(inst0_O[2]), .O(inst3_O));
LUT2 #(.INIT(4'h2)) inst4 (.I0(I[3]), .I1(inst0_O[3]), .O(inst4_O));
LUT2 #(.INIT(4'h2)) inst5 (.I0(I[4]), .I1(inst0_O[4]), .O(inst5_O));
LUT2 #(.INIT(4'h2)) inst6 (.I0(I[5]), .I1(inst0_O[5]), .O(inst6_O));
LUT2 #(.INIT(4'h2)) inst7 (.I0(I[6]), .I1(inst0_O[6]), .O(inst7_O));
LUT2 #(.INIT(4'h2)) inst8 (.I0(I[7]), .I1(inst0_O[7]), .O(inst8_O));
assign O = {inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O};
endmodule

module Encoder8 (input [7:0] I, output [2:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
LUT4 #(.INIT(16'hFFFE)) inst0 (.I0(I[1]), .I1(I[3]), .I2(I[5]), .I3(I[7]), .O(inst0_O));
LUT4 #(.INIT(16'hFFFE)) inst1 (.I0(I[2]), .I1(I[3]), .I2(I[6]), .I3(I[7]), .O(inst1_O));
LUT4 #(.INIT(16'hFFFE)) inst2 (.I0(I[4]), .I1(I[5]), .I2(I[6]), .I3(I[7]), .O(inst2_O));
assign O = {inst2_O,inst1_O,inst0_O};
endmodule

module main (output [2:0] LED, input [7:0] SWITCH);
wire [7:0] inst0_O;
wire [2:0] inst1_O;
Arbiter8 inst0 (.I(SWITCH), .O(inst0_O));
Encoder8 inst1 (.I(inst0_O), .O(inst1_O));
assign LED = inst1_O;
endmodule

