module coreir_reg_arst #(parameter width = 1, parameter arst_posedge = 1, parameter clk_posedge = 1, parameter init = 1) (input clk, input arst, input [width-1:0] in, output [width-1:0] out);
  reg [width-1:0] outReg;
  wire real_rst;
  assign real_rst = arst_posedge ? arst : ~arst;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk, posedge real_rst) begin
    if (real_rst) outReg <= init;
    else outReg <= in;
  end
  assign out = outReg;
endmodule

module test (input ASYNCRESETN, input CLK, input [0:0] In0, output [0:0] Out0, input clk);
wire [0:0] reg_PR_inst0_out;
coreir_reg_arst #(.arst_posedge(0), .clk_posedge(1), .init(1'h0), .width(1)) reg_PR_inst0(.arst(ASYNCRESETN), .clk(clk), .in(In0), .out(reg_PR_inst0_out));
assign Out0 = reg_PR_inst0_out;
endmodule

