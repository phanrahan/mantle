module Decode998 (
    input [7:0] I,
    output O
);
assign O = I == 8'h63;
endmodule

module Decode988 (
    input [7:0] I,
    output O
);
assign O = I == 8'h62;
endmodule

module Decode98 (
    input [7:0] I,
    output O
);
assign O = I == 8'h09;
endmodule

module Decode978 (
    input [7:0] I,
    output O
);
assign O = I == 8'h61;
endmodule

module Decode968 (
    input [7:0] I,
    output O
);
assign O = I == 8'h60;
endmodule

module Decode958 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5f;
endmodule

module Decode948 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5e;
endmodule

module Decode938 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5d;
endmodule

module Decode928 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5c;
endmodule

module Decode918 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5b;
endmodule

module Decode908 (
    input [7:0] I,
    output O
);
assign O = I == 8'h5a;
endmodule

module Decode898 (
    input [7:0] I,
    output O
);
assign O = I == 8'h59;
endmodule

module Decode888 (
    input [7:0] I,
    output O
);
assign O = I == 8'h58;
endmodule

module Decode88 (
    input [7:0] I,
    output O
);
assign O = I == 8'h08;
endmodule

module Decode878 (
    input [7:0] I,
    output O
);
assign O = I == 8'h57;
endmodule

module Decode868 (
    input [7:0] I,
    output O
);
assign O = I == 8'h56;
endmodule

module Decode858 (
    input [7:0] I,
    output O
);
assign O = I == 8'h55;
endmodule

module Decode848 (
    input [7:0] I,
    output O
);
assign O = I == 8'h54;
endmodule

module Decode838 (
    input [7:0] I,
    output O
);
assign O = I == 8'h53;
endmodule

module Decode828 (
    input [7:0] I,
    output O
);
assign O = I == 8'h52;
endmodule

module Decode818 (
    input [7:0] I,
    output O
);
assign O = I == 8'h51;
endmodule

module Decode808 (
    input [7:0] I,
    output O
);
assign O = I == 8'h50;
endmodule

module Decode798 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4f;
endmodule

module Decode788 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4e;
endmodule

module Decode78 (
    input [7:0] I,
    output O
);
assign O = I == 8'h07;
endmodule

module Decode778 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4d;
endmodule

module Decode768 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4c;
endmodule

module Decode758 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4b;
endmodule

module Decode748 (
    input [7:0] I,
    output O
);
assign O = I == 8'h4a;
endmodule

module Decode738 (
    input [7:0] I,
    output O
);
assign O = I == 8'h49;
endmodule

module Decode728 (
    input [7:0] I,
    output O
);
assign O = I == 8'h48;
endmodule

module Decode718 (
    input [7:0] I,
    output O
);
assign O = I == 8'h47;
endmodule

module Decode708 (
    input [7:0] I,
    output O
);
assign O = I == 8'h46;
endmodule

module Decode698 (
    input [7:0] I,
    output O
);
assign O = I == 8'h45;
endmodule

module Decode688 (
    input [7:0] I,
    output O
);
assign O = I == 8'h44;
endmodule

module Decode68 (
    input [7:0] I,
    output O
);
assign O = I == 8'h06;
endmodule

module Decode678 (
    input [7:0] I,
    output O
);
assign O = I == 8'h43;
endmodule

module Decode668 (
    input [7:0] I,
    output O
);
assign O = I == 8'h42;
endmodule

module Decode658 (
    input [7:0] I,
    output O
);
assign O = I == 8'h41;
endmodule

module Decode648 (
    input [7:0] I,
    output O
);
assign O = I == 8'h40;
endmodule

module Decode638 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3f;
endmodule

module Decode628 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3e;
endmodule

module Decode618 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3d;
endmodule

module Decode608 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3c;
endmodule

module Decode598 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3b;
endmodule

module Decode588 (
    input [7:0] I,
    output O
);
assign O = I == 8'h3a;
endmodule

module Decode58 (
    input [7:0] I,
    output O
);
assign O = I == 8'h05;
endmodule

module Decode578 (
    input [7:0] I,
    output O
);
assign O = I == 8'h39;
endmodule

module Decode568 (
    input [7:0] I,
    output O
);
assign O = I == 8'h38;
endmodule

module Decode558 (
    input [7:0] I,
    output O
);
assign O = I == 8'h37;
endmodule

module Decode548 (
    input [7:0] I,
    output O
);
assign O = I == 8'h36;
endmodule

module Decode538 (
    input [7:0] I,
    output O
);
assign O = I == 8'h35;
endmodule

module Decode528 (
    input [7:0] I,
    output O
);
assign O = I == 8'h34;
endmodule

module Decode518 (
    input [7:0] I,
    output O
);
assign O = I == 8'h33;
endmodule

module Decode508 (
    input [7:0] I,
    output O
);
assign O = I == 8'h32;
endmodule

module Decode498 (
    input [7:0] I,
    output O
);
assign O = I == 8'h31;
endmodule

module Decode488 (
    input [7:0] I,
    output O
);
assign O = I == 8'h30;
endmodule

module Decode48 (
    input [7:0] I,
    output O
);
assign O = I == 8'h04;
endmodule

module Decode478 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2f;
endmodule

module Decode468 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2e;
endmodule

module Decode458 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2d;
endmodule

module Decode448 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2c;
endmodule

module Decode438 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2b;
endmodule

module Decode428 (
    input [7:0] I,
    output O
);
assign O = I == 8'h2a;
endmodule

module Decode418 (
    input [7:0] I,
    output O
);
assign O = I == 8'h29;
endmodule

module Decode408 (
    input [7:0] I,
    output O
);
assign O = I == 8'h28;
endmodule

module Decode398 (
    input [7:0] I,
    output O
);
assign O = I == 8'h27;
endmodule

module Decode388 (
    input [7:0] I,
    output O
);
assign O = I == 8'h26;
endmodule

module Decode38 (
    input [7:0] I,
    output O
);
assign O = I == 8'h03;
endmodule

module Decode378 (
    input [7:0] I,
    output O
);
assign O = I == 8'h25;
endmodule

module Decode368 (
    input [7:0] I,
    output O
);
assign O = I == 8'h24;
endmodule

module Decode358 (
    input [7:0] I,
    output O
);
assign O = I == 8'h23;
endmodule

module Decode348 (
    input [7:0] I,
    output O
);
assign O = I == 8'h22;
endmodule

module Decode338 (
    input [7:0] I,
    output O
);
assign O = I == 8'h21;
endmodule

module Decode328 (
    input [7:0] I,
    output O
);
assign O = I == 8'h20;
endmodule

module Decode318 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1f;
endmodule

module Decode308 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1e;
endmodule

module Decode298 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1d;
endmodule

module Decode288 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1c;
endmodule

module Decode28 (
    input [7:0] I,
    output O
);
assign O = I == 8'h02;
endmodule

module Decode278 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1b;
endmodule

module Decode268 (
    input [7:0] I,
    output O
);
assign O = I == 8'h1a;
endmodule

module Decode258 (
    input [7:0] I,
    output O
);
assign O = I == 8'h19;
endmodule

module Decode2558 (
    input [7:0] I,
    output O
);
assign O = I == 8'hff;
endmodule

module Decode2548 (
    input [7:0] I,
    output O
);
assign O = I == 8'hfe;
endmodule

module Decode2538 (
    input [7:0] I,
    output O
);
assign O = I == 8'hfd;
endmodule

module Decode2528 (
    input [7:0] I,
    output O
);
assign O = I == 8'hfc;
endmodule

module Decode2518 (
    input [7:0] I,
    output O
);
assign O = I == 8'hfb;
endmodule

module Decode2508 (
    input [7:0] I,
    output O
);
assign O = I == 8'hfa;
endmodule

module Decode2498 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf9;
endmodule

module Decode2488 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf8;
endmodule

module Decode248 (
    input [7:0] I,
    output O
);
assign O = I == 8'h18;
endmodule

module Decode2478 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf7;
endmodule

module Decode2468 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf6;
endmodule

module Decode2458 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf5;
endmodule

module Decode2448 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf4;
endmodule

module Decode2438 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf3;
endmodule

module Decode2428 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf2;
endmodule

module Decode2418 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf1;
endmodule

module Decode2408 (
    input [7:0] I,
    output O
);
assign O = I == 8'hf0;
endmodule

module Decode2398 (
    input [7:0] I,
    output O
);
assign O = I == 8'hef;
endmodule

module Decode2388 (
    input [7:0] I,
    output O
);
assign O = I == 8'hee;
endmodule

module Decode238 (
    input [7:0] I,
    output O
);
assign O = I == 8'h17;
endmodule

module Decode2378 (
    input [7:0] I,
    output O
);
assign O = I == 8'hed;
endmodule

module Decode2368 (
    input [7:0] I,
    output O
);
assign O = I == 8'hec;
endmodule

module Decode2358 (
    input [7:0] I,
    output O
);
assign O = I == 8'heb;
endmodule

module Decode2348 (
    input [7:0] I,
    output O
);
assign O = I == 8'hea;
endmodule

module Decode2338 (
    input [7:0] I,
    output O
);
assign O = I == 8'he9;
endmodule

module Decode2328 (
    input [7:0] I,
    output O
);
assign O = I == 8'he8;
endmodule

module Decode2318 (
    input [7:0] I,
    output O
);
assign O = I == 8'he7;
endmodule

module Decode2308 (
    input [7:0] I,
    output O
);
assign O = I == 8'he6;
endmodule

module Decode2298 (
    input [7:0] I,
    output O
);
assign O = I == 8'he5;
endmodule

module Decode2288 (
    input [7:0] I,
    output O
);
assign O = I == 8'he4;
endmodule

module Decode228 (
    input [7:0] I,
    output O
);
assign O = I == 8'h16;
endmodule

module Decode2278 (
    input [7:0] I,
    output O
);
assign O = I == 8'he3;
endmodule

module Decode2268 (
    input [7:0] I,
    output O
);
assign O = I == 8'he2;
endmodule

module Decode2258 (
    input [7:0] I,
    output O
);
assign O = I == 8'he1;
endmodule

module Decode2248 (
    input [7:0] I,
    output O
);
assign O = I == 8'he0;
endmodule

module Decode2238 (
    input [7:0] I,
    output O
);
assign O = I == 8'hdf;
endmodule

module Decode2228 (
    input [7:0] I,
    output O
);
assign O = I == 8'hde;
endmodule

module Decode2218 (
    input [7:0] I,
    output O
);
assign O = I == 8'hdd;
endmodule

module Decode2208 (
    input [7:0] I,
    output O
);
assign O = I == 8'hdc;
endmodule

module Decode2198 (
    input [7:0] I,
    output O
);
assign O = I == 8'hdb;
endmodule

module Decode2188 (
    input [7:0] I,
    output O
);
assign O = I == 8'hda;
endmodule

module Decode218 (
    input [7:0] I,
    output O
);
assign O = I == 8'h15;
endmodule

module Decode2178 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd9;
endmodule

module Decode2168 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd8;
endmodule

module Decode2158 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd7;
endmodule

module Decode2148 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd6;
endmodule

module Decode2138 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd5;
endmodule

module Decode2128 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd4;
endmodule

module Decode2118 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd3;
endmodule

module Decode2108 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd2;
endmodule

module Decode2098 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd1;
endmodule

module Decode2088 (
    input [7:0] I,
    output O
);
assign O = I == 8'hd0;
endmodule

module Decode208 (
    input [7:0] I,
    output O
);
assign O = I == 8'h14;
endmodule

module Decode2078 (
    input [7:0] I,
    output O
);
assign O = I == 8'hcf;
endmodule

module Decode2068 (
    input [7:0] I,
    output O
);
assign O = I == 8'hce;
endmodule

module Decode2058 (
    input [7:0] I,
    output O
);
assign O = I == 8'hcd;
endmodule

module Decode2048 (
    input [7:0] I,
    output O
);
assign O = I == 8'hcc;
endmodule

module Decode2038 (
    input [7:0] I,
    output O
);
assign O = I == 8'hcb;
endmodule

module Decode2028 (
    input [7:0] I,
    output O
);
assign O = I == 8'hca;
endmodule

module Decode2018 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc9;
endmodule

module Decode2008 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc8;
endmodule

module Decode1998 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc7;
endmodule

module Decode1988 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc6;
endmodule

module Decode198 (
    input [7:0] I,
    output O
);
assign O = I == 8'h13;
endmodule

module Decode1978 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc5;
endmodule

module Decode1968 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc4;
endmodule

module Decode1958 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc3;
endmodule

module Decode1948 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc2;
endmodule

module Decode1938 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc1;
endmodule

module Decode1928 (
    input [7:0] I,
    output O
);
assign O = I == 8'hc0;
endmodule

module Decode1918 (
    input [7:0] I,
    output O
);
assign O = I == 8'hbf;
endmodule

module Decode1908 (
    input [7:0] I,
    output O
);
assign O = I == 8'hbe;
endmodule

module Decode1898 (
    input [7:0] I,
    output O
);
assign O = I == 8'hbd;
endmodule

module Decode1888 (
    input [7:0] I,
    output O
);
assign O = I == 8'hbc;
endmodule

module Decode188 (
    input [7:0] I,
    output O
);
assign O = I == 8'h12;
endmodule

module Decode1878 (
    input [7:0] I,
    output O
);
assign O = I == 8'hbb;
endmodule

module Decode1868 (
    input [7:0] I,
    output O
);
assign O = I == 8'hba;
endmodule

module Decode1858 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb9;
endmodule

module Decode1848 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb8;
endmodule

module Decode1838 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb7;
endmodule

module Decode1828 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb6;
endmodule

module Decode1818 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb5;
endmodule

module Decode1808 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb4;
endmodule

module Decode18 (
    input [7:0] I,
    output O
);
assign O = I == 8'h01;
endmodule

module Decode1798 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb3;
endmodule

module Decode1788 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb2;
endmodule

module Decode178 (
    input [7:0] I,
    output O
);
assign O = I == 8'h11;
endmodule

module Decode1778 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb1;
endmodule

module Decode1768 (
    input [7:0] I,
    output O
);
assign O = I == 8'hb0;
endmodule

module Decode1758 (
    input [7:0] I,
    output O
);
assign O = I == 8'haf;
endmodule

module Decode1748 (
    input [7:0] I,
    output O
);
assign O = I == 8'hae;
endmodule

module Decode1738 (
    input [7:0] I,
    output O
);
assign O = I == 8'had;
endmodule

module Decode1728 (
    input [7:0] I,
    output O
);
assign O = I == 8'hac;
endmodule

module Decode1718 (
    input [7:0] I,
    output O
);
assign O = I == 8'hab;
endmodule

module Decode1708 (
    input [7:0] I,
    output O
);
assign O = I == 8'haa;
endmodule

module Decode1698 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha9;
endmodule

module Decode1688 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha8;
endmodule

module Decode168 (
    input [7:0] I,
    output O
);
assign O = I == 8'h10;
endmodule

module Decode1678 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha7;
endmodule

module Decode1668 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha6;
endmodule

module Decode1658 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha5;
endmodule

module Decode1648 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha4;
endmodule

module Decode1638 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha3;
endmodule

module Decode1628 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha2;
endmodule

module Decode1618 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha1;
endmodule

module Decode1608 (
    input [7:0] I,
    output O
);
assign O = I == 8'ha0;
endmodule

module Decode1598 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9f;
endmodule

module Decode1588 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9e;
endmodule

module Decode158 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0f;
endmodule

module Decode1578 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9d;
endmodule

module Decode1568 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9c;
endmodule

module Decode1558 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9b;
endmodule

module Decode1548 (
    input [7:0] I,
    output O
);
assign O = I == 8'h9a;
endmodule

module Decode1538 (
    input [7:0] I,
    output O
);
assign O = I == 8'h99;
endmodule

module Decode1528 (
    input [7:0] I,
    output O
);
assign O = I == 8'h98;
endmodule

module Decode1518 (
    input [7:0] I,
    output O
);
assign O = I == 8'h97;
endmodule

module Decode1508 (
    input [7:0] I,
    output O
);
assign O = I == 8'h96;
endmodule

module Decode1498 (
    input [7:0] I,
    output O
);
assign O = I == 8'h95;
endmodule

module Decode1488 (
    input [7:0] I,
    output O
);
assign O = I == 8'h94;
endmodule

module Decode148 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0e;
endmodule

module Decode1478 (
    input [7:0] I,
    output O
);
assign O = I == 8'h93;
endmodule

module Decode1468 (
    input [7:0] I,
    output O
);
assign O = I == 8'h92;
endmodule

module Decode1458 (
    input [7:0] I,
    output O
);
assign O = I == 8'h91;
endmodule

module Decode1448 (
    input [7:0] I,
    output O
);
assign O = I == 8'h90;
endmodule

module Decode1438 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8f;
endmodule

module Decode1428 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8e;
endmodule

module Decode1418 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8d;
endmodule

module Decode1408 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8c;
endmodule

module Decode1398 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8b;
endmodule

module Decode1388 (
    input [7:0] I,
    output O
);
assign O = I == 8'h8a;
endmodule

module Decode138 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0d;
endmodule

module Decode1378 (
    input [7:0] I,
    output O
);
assign O = I == 8'h89;
endmodule

module Decode1368 (
    input [7:0] I,
    output O
);
assign O = I == 8'h88;
endmodule

module Decode1358 (
    input [7:0] I,
    output O
);
assign O = I == 8'h87;
endmodule

module Decode1348 (
    input [7:0] I,
    output O
);
assign O = I == 8'h86;
endmodule

module Decode1338 (
    input [7:0] I,
    output O
);
assign O = I == 8'h85;
endmodule

module Decode1328 (
    input [7:0] I,
    output O
);
assign O = I == 8'h84;
endmodule

module Decode1318 (
    input [7:0] I,
    output O
);
assign O = I == 8'h83;
endmodule

module Decode1308 (
    input [7:0] I,
    output O
);
assign O = I == 8'h82;
endmodule

module Decode1298 (
    input [7:0] I,
    output O
);
assign O = I == 8'h81;
endmodule

module Decode1288 (
    input [7:0] I,
    output O
);
assign O = I == 8'h80;
endmodule

module Decode128 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0c;
endmodule

module Decode1278 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7f;
endmodule

module Decode1268 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7e;
endmodule

module Decode1258 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7d;
endmodule

module Decode1248 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7c;
endmodule

module Decode1238 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7b;
endmodule

module Decode1228 (
    input [7:0] I,
    output O
);
assign O = I == 8'h7a;
endmodule

module Decode1218 (
    input [7:0] I,
    output O
);
assign O = I == 8'h79;
endmodule

module Decode1208 (
    input [7:0] I,
    output O
);
assign O = I == 8'h78;
endmodule

module Decode1198 (
    input [7:0] I,
    output O
);
assign O = I == 8'h77;
endmodule

module Decode1188 (
    input [7:0] I,
    output O
);
assign O = I == 8'h76;
endmodule

module Decode118 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0b;
endmodule

module Decode1178 (
    input [7:0] I,
    output O
);
assign O = I == 8'h75;
endmodule

module Decode1168 (
    input [7:0] I,
    output O
);
assign O = I == 8'h74;
endmodule

module Decode1158 (
    input [7:0] I,
    output O
);
assign O = I == 8'h73;
endmodule

module Decode1148 (
    input [7:0] I,
    output O
);
assign O = I == 8'h72;
endmodule

module Decode1138 (
    input [7:0] I,
    output O
);
assign O = I == 8'h71;
endmodule

module Decode1128 (
    input [7:0] I,
    output O
);
assign O = I == 8'h70;
endmodule

module Decode1118 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6f;
endmodule

module Decode1108 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6e;
endmodule

module Decode1098 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6d;
endmodule

module Decode1088 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6c;
endmodule

module Decode108 (
    input [7:0] I,
    output O
);
assign O = I == 8'h0a;
endmodule

module Decode1078 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6b;
endmodule

module Decode1068 (
    input [7:0] I,
    output O
);
assign O = I == 8'h6a;
endmodule

module Decode1058 (
    input [7:0] I,
    output O
);
assign O = I == 8'h69;
endmodule

module Decode1048 (
    input [7:0] I,
    output O
);
assign O = I == 8'h68;
endmodule

module Decode1038 (
    input [7:0] I,
    output O
);
assign O = I == 8'h67;
endmodule

module Decode1028 (
    input [7:0] I,
    output O
);
assign O = I == 8'h66;
endmodule

module Decode1018 (
    input [7:0] I,
    output O
);
assign O = I == 8'h65;
endmodule

module Decode1008 (
    input [7:0] I,
    output O
);
assign O = I == 8'h64;
endmodule

module Decode08 (
    input [7:0] I,
    output O
);
assign O = I == 8'h00;
endmodule

module Decoder8 (
    input [7:0] I,
    output [255:0] O
);
wire [7:0] Decode08_inst0_I;
wire Decode08_inst0_O;
wire [7:0] Decode1008_inst0_I;
wire Decode1008_inst0_O;
wire [7:0] Decode1018_inst0_I;
wire Decode1018_inst0_O;
wire [7:0] Decode1028_inst0_I;
wire Decode1028_inst0_O;
wire [7:0] Decode1038_inst0_I;
wire Decode1038_inst0_O;
wire [7:0] Decode1048_inst0_I;
wire Decode1048_inst0_O;
wire [7:0] Decode1058_inst0_I;
wire Decode1058_inst0_O;
wire [7:0] Decode1068_inst0_I;
wire Decode1068_inst0_O;
wire [7:0] Decode1078_inst0_I;
wire Decode1078_inst0_O;
wire [7:0] Decode1088_inst0_I;
wire Decode1088_inst0_O;
wire [7:0] Decode108_inst0_I;
wire Decode108_inst0_O;
wire [7:0] Decode1098_inst0_I;
wire Decode1098_inst0_O;
wire [7:0] Decode1108_inst0_I;
wire Decode1108_inst0_O;
wire [7:0] Decode1118_inst0_I;
wire Decode1118_inst0_O;
wire [7:0] Decode1128_inst0_I;
wire Decode1128_inst0_O;
wire [7:0] Decode1138_inst0_I;
wire Decode1138_inst0_O;
wire [7:0] Decode1148_inst0_I;
wire Decode1148_inst0_O;
wire [7:0] Decode1158_inst0_I;
wire Decode1158_inst0_O;
wire [7:0] Decode1168_inst0_I;
wire Decode1168_inst0_O;
wire [7:0] Decode1178_inst0_I;
wire Decode1178_inst0_O;
wire [7:0] Decode1188_inst0_I;
wire Decode1188_inst0_O;
wire [7:0] Decode118_inst0_I;
wire Decode118_inst0_O;
wire [7:0] Decode1198_inst0_I;
wire Decode1198_inst0_O;
wire [7:0] Decode1208_inst0_I;
wire Decode1208_inst0_O;
wire [7:0] Decode1218_inst0_I;
wire Decode1218_inst0_O;
wire [7:0] Decode1228_inst0_I;
wire Decode1228_inst0_O;
wire [7:0] Decode1238_inst0_I;
wire Decode1238_inst0_O;
wire [7:0] Decode1248_inst0_I;
wire Decode1248_inst0_O;
wire [7:0] Decode1258_inst0_I;
wire Decode1258_inst0_O;
wire [7:0] Decode1268_inst0_I;
wire Decode1268_inst0_O;
wire [7:0] Decode1278_inst0_I;
wire Decode1278_inst0_O;
wire [7:0] Decode1288_inst0_I;
wire Decode1288_inst0_O;
wire [7:0] Decode128_inst0_I;
wire Decode128_inst0_O;
wire [7:0] Decode1298_inst0_I;
wire Decode1298_inst0_O;
wire [7:0] Decode1308_inst0_I;
wire Decode1308_inst0_O;
wire [7:0] Decode1318_inst0_I;
wire Decode1318_inst0_O;
wire [7:0] Decode1328_inst0_I;
wire Decode1328_inst0_O;
wire [7:0] Decode1338_inst0_I;
wire Decode1338_inst0_O;
wire [7:0] Decode1348_inst0_I;
wire Decode1348_inst0_O;
wire [7:0] Decode1358_inst0_I;
wire Decode1358_inst0_O;
wire [7:0] Decode1368_inst0_I;
wire Decode1368_inst0_O;
wire [7:0] Decode1378_inst0_I;
wire Decode1378_inst0_O;
wire [7:0] Decode1388_inst0_I;
wire Decode1388_inst0_O;
wire [7:0] Decode138_inst0_I;
wire Decode138_inst0_O;
wire [7:0] Decode1398_inst0_I;
wire Decode1398_inst0_O;
wire [7:0] Decode1408_inst0_I;
wire Decode1408_inst0_O;
wire [7:0] Decode1418_inst0_I;
wire Decode1418_inst0_O;
wire [7:0] Decode1428_inst0_I;
wire Decode1428_inst0_O;
wire [7:0] Decode1438_inst0_I;
wire Decode1438_inst0_O;
wire [7:0] Decode1448_inst0_I;
wire Decode1448_inst0_O;
wire [7:0] Decode1458_inst0_I;
wire Decode1458_inst0_O;
wire [7:0] Decode1468_inst0_I;
wire Decode1468_inst0_O;
wire [7:0] Decode1478_inst0_I;
wire Decode1478_inst0_O;
wire [7:0] Decode1488_inst0_I;
wire Decode1488_inst0_O;
wire [7:0] Decode148_inst0_I;
wire Decode148_inst0_O;
wire [7:0] Decode1498_inst0_I;
wire Decode1498_inst0_O;
wire [7:0] Decode1508_inst0_I;
wire Decode1508_inst0_O;
wire [7:0] Decode1518_inst0_I;
wire Decode1518_inst0_O;
wire [7:0] Decode1528_inst0_I;
wire Decode1528_inst0_O;
wire [7:0] Decode1538_inst0_I;
wire Decode1538_inst0_O;
wire [7:0] Decode1548_inst0_I;
wire Decode1548_inst0_O;
wire [7:0] Decode1558_inst0_I;
wire Decode1558_inst0_O;
wire [7:0] Decode1568_inst0_I;
wire Decode1568_inst0_O;
wire [7:0] Decode1578_inst0_I;
wire Decode1578_inst0_O;
wire [7:0] Decode1588_inst0_I;
wire Decode1588_inst0_O;
wire [7:0] Decode158_inst0_I;
wire Decode158_inst0_O;
wire [7:0] Decode1598_inst0_I;
wire Decode1598_inst0_O;
wire [7:0] Decode1608_inst0_I;
wire Decode1608_inst0_O;
wire [7:0] Decode1618_inst0_I;
wire Decode1618_inst0_O;
wire [7:0] Decode1628_inst0_I;
wire Decode1628_inst0_O;
wire [7:0] Decode1638_inst0_I;
wire Decode1638_inst0_O;
wire [7:0] Decode1648_inst0_I;
wire Decode1648_inst0_O;
wire [7:0] Decode1658_inst0_I;
wire Decode1658_inst0_O;
wire [7:0] Decode1668_inst0_I;
wire Decode1668_inst0_O;
wire [7:0] Decode1678_inst0_I;
wire Decode1678_inst0_O;
wire [7:0] Decode1688_inst0_I;
wire Decode1688_inst0_O;
wire [7:0] Decode168_inst0_I;
wire Decode168_inst0_O;
wire [7:0] Decode1698_inst0_I;
wire Decode1698_inst0_O;
wire [7:0] Decode1708_inst0_I;
wire Decode1708_inst0_O;
wire [7:0] Decode1718_inst0_I;
wire Decode1718_inst0_O;
wire [7:0] Decode1728_inst0_I;
wire Decode1728_inst0_O;
wire [7:0] Decode1738_inst0_I;
wire Decode1738_inst0_O;
wire [7:0] Decode1748_inst0_I;
wire Decode1748_inst0_O;
wire [7:0] Decode1758_inst0_I;
wire Decode1758_inst0_O;
wire [7:0] Decode1768_inst0_I;
wire Decode1768_inst0_O;
wire [7:0] Decode1778_inst0_I;
wire Decode1778_inst0_O;
wire [7:0] Decode1788_inst0_I;
wire Decode1788_inst0_O;
wire [7:0] Decode178_inst0_I;
wire Decode178_inst0_O;
wire [7:0] Decode1798_inst0_I;
wire Decode1798_inst0_O;
wire [7:0] Decode1808_inst0_I;
wire Decode1808_inst0_O;
wire [7:0] Decode1818_inst0_I;
wire Decode1818_inst0_O;
wire [7:0] Decode1828_inst0_I;
wire Decode1828_inst0_O;
wire [7:0] Decode1838_inst0_I;
wire Decode1838_inst0_O;
wire [7:0] Decode1848_inst0_I;
wire Decode1848_inst0_O;
wire [7:0] Decode1858_inst0_I;
wire Decode1858_inst0_O;
wire [7:0] Decode1868_inst0_I;
wire Decode1868_inst0_O;
wire [7:0] Decode1878_inst0_I;
wire Decode1878_inst0_O;
wire [7:0] Decode1888_inst0_I;
wire Decode1888_inst0_O;
wire [7:0] Decode188_inst0_I;
wire Decode188_inst0_O;
wire [7:0] Decode1898_inst0_I;
wire Decode1898_inst0_O;
wire [7:0] Decode18_inst0_I;
wire Decode18_inst0_O;
wire [7:0] Decode1908_inst0_I;
wire Decode1908_inst0_O;
wire [7:0] Decode1918_inst0_I;
wire Decode1918_inst0_O;
wire [7:0] Decode1928_inst0_I;
wire Decode1928_inst0_O;
wire [7:0] Decode1938_inst0_I;
wire Decode1938_inst0_O;
wire [7:0] Decode1948_inst0_I;
wire Decode1948_inst0_O;
wire [7:0] Decode1958_inst0_I;
wire Decode1958_inst0_O;
wire [7:0] Decode1968_inst0_I;
wire Decode1968_inst0_O;
wire [7:0] Decode1978_inst0_I;
wire Decode1978_inst0_O;
wire [7:0] Decode1988_inst0_I;
wire Decode1988_inst0_O;
wire [7:0] Decode198_inst0_I;
wire Decode198_inst0_O;
wire [7:0] Decode1998_inst0_I;
wire Decode1998_inst0_O;
wire [7:0] Decode2008_inst0_I;
wire Decode2008_inst0_O;
wire [7:0] Decode2018_inst0_I;
wire Decode2018_inst0_O;
wire [7:0] Decode2028_inst0_I;
wire Decode2028_inst0_O;
wire [7:0] Decode2038_inst0_I;
wire Decode2038_inst0_O;
wire [7:0] Decode2048_inst0_I;
wire Decode2048_inst0_O;
wire [7:0] Decode2058_inst0_I;
wire Decode2058_inst0_O;
wire [7:0] Decode2068_inst0_I;
wire Decode2068_inst0_O;
wire [7:0] Decode2078_inst0_I;
wire Decode2078_inst0_O;
wire [7:0] Decode2088_inst0_I;
wire Decode2088_inst0_O;
wire [7:0] Decode208_inst0_I;
wire Decode208_inst0_O;
wire [7:0] Decode2098_inst0_I;
wire Decode2098_inst0_O;
wire [7:0] Decode2108_inst0_I;
wire Decode2108_inst0_O;
wire [7:0] Decode2118_inst0_I;
wire Decode2118_inst0_O;
wire [7:0] Decode2128_inst0_I;
wire Decode2128_inst0_O;
wire [7:0] Decode2138_inst0_I;
wire Decode2138_inst0_O;
wire [7:0] Decode2148_inst0_I;
wire Decode2148_inst0_O;
wire [7:0] Decode2158_inst0_I;
wire Decode2158_inst0_O;
wire [7:0] Decode2168_inst0_I;
wire Decode2168_inst0_O;
wire [7:0] Decode2178_inst0_I;
wire Decode2178_inst0_O;
wire [7:0] Decode2188_inst0_I;
wire Decode2188_inst0_O;
wire [7:0] Decode218_inst0_I;
wire Decode218_inst0_O;
wire [7:0] Decode2198_inst0_I;
wire Decode2198_inst0_O;
wire [7:0] Decode2208_inst0_I;
wire Decode2208_inst0_O;
wire [7:0] Decode2218_inst0_I;
wire Decode2218_inst0_O;
wire [7:0] Decode2228_inst0_I;
wire Decode2228_inst0_O;
wire [7:0] Decode2238_inst0_I;
wire Decode2238_inst0_O;
wire [7:0] Decode2248_inst0_I;
wire Decode2248_inst0_O;
wire [7:0] Decode2258_inst0_I;
wire Decode2258_inst0_O;
wire [7:0] Decode2268_inst0_I;
wire Decode2268_inst0_O;
wire [7:0] Decode2278_inst0_I;
wire Decode2278_inst0_O;
wire [7:0] Decode2288_inst0_I;
wire Decode2288_inst0_O;
wire [7:0] Decode228_inst0_I;
wire Decode228_inst0_O;
wire [7:0] Decode2298_inst0_I;
wire Decode2298_inst0_O;
wire [7:0] Decode2308_inst0_I;
wire Decode2308_inst0_O;
wire [7:0] Decode2318_inst0_I;
wire Decode2318_inst0_O;
wire [7:0] Decode2328_inst0_I;
wire Decode2328_inst0_O;
wire [7:0] Decode2338_inst0_I;
wire Decode2338_inst0_O;
wire [7:0] Decode2348_inst0_I;
wire Decode2348_inst0_O;
wire [7:0] Decode2358_inst0_I;
wire Decode2358_inst0_O;
wire [7:0] Decode2368_inst0_I;
wire Decode2368_inst0_O;
wire [7:0] Decode2378_inst0_I;
wire Decode2378_inst0_O;
wire [7:0] Decode2388_inst0_I;
wire Decode2388_inst0_O;
wire [7:0] Decode238_inst0_I;
wire Decode238_inst0_O;
wire [7:0] Decode2398_inst0_I;
wire Decode2398_inst0_O;
wire [7:0] Decode2408_inst0_I;
wire Decode2408_inst0_O;
wire [7:0] Decode2418_inst0_I;
wire Decode2418_inst0_O;
wire [7:0] Decode2428_inst0_I;
wire Decode2428_inst0_O;
wire [7:0] Decode2438_inst0_I;
wire Decode2438_inst0_O;
wire [7:0] Decode2448_inst0_I;
wire Decode2448_inst0_O;
wire [7:0] Decode2458_inst0_I;
wire Decode2458_inst0_O;
wire [7:0] Decode2468_inst0_I;
wire Decode2468_inst0_O;
wire [7:0] Decode2478_inst0_I;
wire Decode2478_inst0_O;
wire [7:0] Decode2488_inst0_I;
wire Decode2488_inst0_O;
wire [7:0] Decode248_inst0_I;
wire Decode248_inst0_O;
wire [7:0] Decode2498_inst0_I;
wire Decode2498_inst0_O;
wire [7:0] Decode2508_inst0_I;
wire Decode2508_inst0_O;
wire [7:0] Decode2518_inst0_I;
wire Decode2518_inst0_O;
wire [7:0] Decode2528_inst0_I;
wire Decode2528_inst0_O;
wire [7:0] Decode2538_inst0_I;
wire Decode2538_inst0_O;
wire [7:0] Decode2548_inst0_I;
wire Decode2548_inst0_O;
wire [7:0] Decode2558_inst0_I;
wire Decode2558_inst0_O;
wire [7:0] Decode258_inst0_I;
wire Decode258_inst0_O;
wire [7:0] Decode268_inst0_I;
wire Decode268_inst0_O;
wire [7:0] Decode278_inst0_I;
wire Decode278_inst0_O;
wire [7:0] Decode288_inst0_I;
wire Decode288_inst0_O;
wire [7:0] Decode28_inst0_I;
wire Decode28_inst0_O;
wire [7:0] Decode298_inst0_I;
wire Decode298_inst0_O;
wire [7:0] Decode308_inst0_I;
wire Decode308_inst0_O;
wire [7:0] Decode318_inst0_I;
wire Decode318_inst0_O;
wire [7:0] Decode328_inst0_I;
wire Decode328_inst0_O;
wire [7:0] Decode338_inst0_I;
wire Decode338_inst0_O;
wire [7:0] Decode348_inst0_I;
wire Decode348_inst0_O;
wire [7:0] Decode358_inst0_I;
wire Decode358_inst0_O;
wire [7:0] Decode368_inst0_I;
wire Decode368_inst0_O;
wire [7:0] Decode378_inst0_I;
wire Decode378_inst0_O;
wire [7:0] Decode388_inst0_I;
wire Decode388_inst0_O;
wire [7:0] Decode38_inst0_I;
wire Decode38_inst0_O;
wire [7:0] Decode398_inst0_I;
wire Decode398_inst0_O;
wire [7:0] Decode408_inst0_I;
wire Decode408_inst0_O;
wire [7:0] Decode418_inst0_I;
wire Decode418_inst0_O;
wire [7:0] Decode428_inst0_I;
wire Decode428_inst0_O;
wire [7:0] Decode438_inst0_I;
wire Decode438_inst0_O;
wire [7:0] Decode448_inst0_I;
wire Decode448_inst0_O;
wire [7:0] Decode458_inst0_I;
wire Decode458_inst0_O;
wire [7:0] Decode468_inst0_I;
wire Decode468_inst0_O;
wire [7:0] Decode478_inst0_I;
wire Decode478_inst0_O;
wire [7:0] Decode488_inst0_I;
wire Decode488_inst0_O;
wire [7:0] Decode48_inst0_I;
wire Decode48_inst0_O;
wire [7:0] Decode498_inst0_I;
wire Decode498_inst0_O;
wire [7:0] Decode508_inst0_I;
wire Decode508_inst0_O;
wire [7:0] Decode518_inst0_I;
wire Decode518_inst0_O;
wire [7:0] Decode528_inst0_I;
wire Decode528_inst0_O;
wire [7:0] Decode538_inst0_I;
wire Decode538_inst0_O;
wire [7:0] Decode548_inst0_I;
wire Decode548_inst0_O;
wire [7:0] Decode558_inst0_I;
wire Decode558_inst0_O;
wire [7:0] Decode568_inst0_I;
wire Decode568_inst0_O;
wire [7:0] Decode578_inst0_I;
wire Decode578_inst0_O;
wire [7:0] Decode588_inst0_I;
wire Decode588_inst0_O;
wire [7:0] Decode58_inst0_I;
wire Decode58_inst0_O;
wire [7:0] Decode598_inst0_I;
wire Decode598_inst0_O;
wire [7:0] Decode608_inst0_I;
wire Decode608_inst0_O;
wire [7:0] Decode618_inst0_I;
wire Decode618_inst0_O;
wire [7:0] Decode628_inst0_I;
wire Decode628_inst0_O;
wire [7:0] Decode638_inst0_I;
wire Decode638_inst0_O;
wire [7:0] Decode648_inst0_I;
wire Decode648_inst0_O;
wire [7:0] Decode658_inst0_I;
wire Decode658_inst0_O;
wire [7:0] Decode668_inst0_I;
wire Decode668_inst0_O;
wire [7:0] Decode678_inst0_I;
wire Decode678_inst0_O;
wire [7:0] Decode688_inst0_I;
wire Decode688_inst0_O;
wire [7:0] Decode68_inst0_I;
wire Decode68_inst0_O;
wire [7:0] Decode698_inst0_I;
wire Decode698_inst0_O;
wire [7:0] Decode708_inst0_I;
wire Decode708_inst0_O;
wire [7:0] Decode718_inst0_I;
wire Decode718_inst0_O;
wire [7:0] Decode728_inst0_I;
wire Decode728_inst0_O;
wire [7:0] Decode738_inst0_I;
wire Decode738_inst0_O;
wire [7:0] Decode748_inst0_I;
wire Decode748_inst0_O;
wire [7:0] Decode758_inst0_I;
wire Decode758_inst0_O;
wire [7:0] Decode768_inst0_I;
wire Decode768_inst0_O;
wire [7:0] Decode778_inst0_I;
wire Decode778_inst0_O;
wire [7:0] Decode788_inst0_I;
wire Decode788_inst0_O;
wire [7:0] Decode78_inst0_I;
wire Decode78_inst0_O;
wire [7:0] Decode798_inst0_I;
wire Decode798_inst0_O;
wire [7:0] Decode808_inst0_I;
wire Decode808_inst0_O;
wire [7:0] Decode818_inst0_I;
wire Decode818_inst0_O;
wire [7:0] Decode828_inst0_I;
wire Decode828_inst0_O;
wire [7:0] Decode838_inst0_I;
wire Decode838_inst0_O;
wire [7:0] Decode848_inst0_I;
wire Decode848_inst0_O;
wire [7:0] Decode858_inst0_I;
wire Decode858_inst0_O;
wire [7:0] Decode868_inst0_I;
wire Decode868_inst0_O;
wire [7:0] Decode878_inst0_I;
wire Decode878_inst0_O;
wire [7:0] Decode888_inst0_I;
wire Decode888_inst0_O;
wire [7:0] Decode88_inst0_I;
wire Decode88_inst0_O;
wire [7:0] Decode898_inst0_I;
wire Decode898_inst0_O;
wire [7:0] Decode908_inst0_I;
wire Decode908_inst0_O;
wire [7:0] Decode918_inst0_I;
wire Decode918_inst0_O;
wire [7:0] Decode928_inst0_I;
wire Decode928_inst0_O;
wire [7:0] Decode938_inst0_I;
wire Decode938_inst0_O;
wire [7:0] Decode948_inst0_I;
wire Decode948_inst0_O;
wire [7:0] Decode958_inst0_I;
wire Decode958_inst0_O;
wire [7:0] Decode968_inst0_I;
wire Decode968_inst0_O;
wire [7:0] Decode978_inst0_I;
wire Decode978_inst0_O;
wire [7:0] Decode988_inst0_I;
wire Decode988_inst0_O;
wire [7:0] Decode98_inst0_I;
wire Decode98_inst0_O;
wire [7:0] Decode998_inst0_I;
wire Decode998_inst0_O;
assign Decode08_inst0_I = I;
Decode08 Decode08_inst0 (
    .I(Decode08_inst0_I),
    .O(Decode08_inst0_O)
);
assign Decode1008_inst0_I = I;
Decode1008 Decode1008_inst0 (
    .I(Decode1008_inst0_I),
    .O(Decode1008_inst0_O)
);
assign Decode1018_inst0_I = I;
Decode1018 Decode1018_inst0 (
    .I(Decode1018_inst0_I),
    .O(Decode1018_inst0_O)
);
assign Decode1028_inst0_I = I;
Decode1028 Decode1028_inst0 (
    .I(Decode1028_inst0_I),
    .O(Decode1028_inst0_O)
);
assign Decode1038_inst0_I = I;
Decode1038 Decode1038_inst0 (
    .I(Decode1038_inst0_I),
    .O(Decode1038_inst0_O)
);
assign Decode1048_inst0_I = I;
Decode1048 Decode1048_inst0 (
    .I(Decode1048_inst0_I),
    .O(Decode1048_inst0_O)
);
assign Decode1058_inst0_I = I;
Decode1058 Decode1058_inst0 (
    .I(Decode1058_inst0_I),
    .O(Decode1058_inst0_O)
);
assign Decode1068_inst0_I = I;
Decode1068 Decode1068_inst0 (
    .I(Decode1068_inst0_I),
    .O(Decode1068_inst0_O)
);
assign Decode1078_inst0_I = I;
Decode1078 Decode1078_inst0 (
    .I(Decode1078_inst0_I),
    .O(Decode1078_inst0_O)
);
assign Decode1088_inst0_I = I;
Decode1088 Decode1088_inst0 (
    .I(Decode1088_inst0_I),
    .O(Decode1088_inst0_O)
);
assign Decode108_inst0_I = I;
Decode108 Decode108_inst0 (
    .I(Decode108_inst0_I),
    .O(Decode108_inst0_O)
);
assign Decode1098_inst0_I = I;
Decode1098 Decode1098_inst0 (
    .I(Decode1098_inst0_I),
    .O(Decode1098_inst0_O)
);
assign Decode1108_inst0_I = I;
Decode1108 Decode1108_inst0 (
    .I(Decode1108_inst0_I),
    .O(Decode1108_inst0_O)
);
assign Decode1118_inst0_I = I;
Decode1118 Decode1118_inst0 (
    .I(Decode1118_inst0_I),
    .O(Decode1118_inst0_O)
);
assign Decode1128_inst0_I = I;
Decode1128 Decode1128_inst0 (
    .I(Decode1128_inst0_I),
    .O(Decode1128_inst0_O)
);
assign Decode1138_inst0_I = I;
Decode1138 Decode1138_inst0 (
    .I(Decode1138_inst0_I),
    .O(Decode1138_inst0_O)
);
assign Decode1148_inst0_I = I;
Decode1148 Decode1148_inst0 (
    .I(Decode1148_inst0_I),
    .O(Decode1148_inst0_O)
);
assign Decode1158_inst0_I = I;
Decode1158 Decode1158_inst0 (
    .I(Decode1158_inst0_I),
    .O(Decode1158_inst0_O)
);
assign Decode1168_inst0_I = I;
Decode1168 Decode1168_inst0 (
    .I(Decode1168_inst0_I),
    .O(Decode1168_inst0_O)
);
assign Decode1178_inst0_I = I;
Decode1178 Decode1178_inst0 (
    .I(Decode1178_inst0_I),
    .O(Decode1178_inst0_O)
);
assign Decode1188_inst0_I = I;
Decode1188 Decode1188_inst0 (
    .I(Decode1188_inst0_I),
    .O(Decode1188_inst0_O)
);
assign Decode118_inst0_I = I;
Decode118 Decode118_inst0 (
    .I(Decode118_inst0_I),
    .O(Decode118_inst0_O)
);
assign Decode1198_inst0_I = I;
Decode1198 Decode1198_inst0 (
    .I(Decode1198_inst0_I),
    .O(Decode1198_inst0_O)
);
assign Decode1208_inst0_I = I;
Decode1208 Decode1208_inst0 (
    .I(Decode1208_inst0_I),
    .O(Decode1208_inst0_O)
);
assign Decode1218_inst0_I = I;
Decode1218 Decode1218_inst0 (
    .I(Decode1218_inst0_I),
    .O(Decode1218_inst0_O)
);
assign Decode1228_inst0_I = I;
Decode1228 Decode1228_inst0 (
    .I(Decode1228_inst0_I),
    .O(Decode1228_inst0_O)
);
assign Decode1238_inst0_I = I;
Decode1238 Decode1238_inst0 (
    .I(Decode1238_inst0_I),
    .O(Decode1238_inst0_O)
);
assign Decode1248_inst0_I = I;
Decode1248 Decode1248_inst0 (
    .I(Decode1248_inst0_I),
    .O(Decode1248_inst0_O)
);
assign Decode1258_inst0_I = I;
Decode1258 Decode1258_inst0 (
    .I(Decode1258_inst0_I),
    .O(Decode1258_inst0_O)
);
assign Decode1268_inst0_I = I;
Decode1268 Decode1268_inst0 (
    .I(Decode1268_inst0_I),
    .O(Decode1268_inst0_O)
);
assign Decode1278_inst0_I = I;
Decode1278 Decode1278_inst0 (
    .I(Decode1278_inst0_I),
    .O(Decode1278_inst0_O)
);
assign Decode1288_inst0_I = I;
Decode1288 Decode1288_inst0 (
    .I(Decode1288_inst0_I),
    .O(Decode1288_inst0_O)
);
assign Decode128_inst0_I = I;
Decode128 Decode128_inst0 (
    .I(Decode128_inst0_I),
    .O(Decode128_inst0_O)
);
assign Decode1298_inst0_I = I;
Decode1298 Decode1298_inst0 (
    .I(Decode1298_inst0_I),
    .O(Decode1298_inst0_O)
);
assign Decode1308_inst0_I = I;
Decode1308 Decode1308_inst0 (
    .I(Decode1308_inst0_I),
    .O(Decode1308_inst0_O)
);
assign Decode1318_inst0_I = I;
Decode1318 Decode1318_inst0 (
    .I(Decode1318_inst0_I),
    .O(Decode1318_inst0_O)
);
assign Decode1328_inst0_I = I;
Decode1328 Decode1328_inst0 (
    .I(Decode1328_inst0_I),
    .O(Decode1328_inst0_O)
);
assign Decode1338_inst0_I = I;
Decode1338 Decode1338_inst0 (
    .I(Decode1338_inst0_I),
    .O(Decode1338_inst0_O)
);
assign Decode1348_inst0_I = I;
Decode1348 Decode1348_inst0 (
    .I(Decode1348_inst0_I),
    .O(Decode1348_inst0_O)
);
assign Decode1358_inst0_I = I;
Decode1358 Decode1358_inst0 (
    .I(Decode1358_inst0_I),
    .O(Decode1358_inst0_O)
);
assign Decode1368_inst0_I = I;
Decode1368 Decode1368_inst0 (
    .I(Decode1368_inst0_I),
    .O(Decode1368_inst0_O)
);
assign Decode1378_inst0_I = I;
Decode1378 Decode1378_inst0 (
    .I(Decode1378_inst0_I),
    .O(Decode1378_inst0_O)
);
assign Decode1388_inst0_I = I;
Decode1388 Decode1388_inst0 (
    .I(Decode1388_inst0_I),
    .O(Decode1388_inst0_O)
);
assign Decode138_inst0_I = I;
Decode138 Decode138_inst0 (
    .I(Decode138_inst0_I),
    .O(Decode138_inst0_O)
);
assign Decode1398_inst0_I = I;
Decode1398 Decode1398_inst0 (
    .I(Decode1398_inst0_I),
    .O(Decode1398_inst0_O)
);
assign Decode1408_inst0_I = I;
Decode1408 Decode1408_inst0 (
    .I(Decode1408_inst0_I),
    .O(Decode1408_inst0_O)
);
assign Decode1418_inst0_I = I;
Decode1418 Decode1418_inst0 (
    .I(Decode1418_inst0_I),
    .O(Decode1418_inst0_O)
);
assign Decode1428_inst0_I = I;
Decode1428 Decode1428_inst0 (
    .I(Decode1428_inst0_I),
    .O(Decode1428_inst0_O)
);
assign Decode1438_inst0_I = I;
Decode1438 Decode1438_inst0 (
    .I(Decode1438_inst0_I),
    .O(Decode1438_inst0_O)
);
assign Decode1448_inst0_I = I;
Decode1448 Decode1448_inst0 (
    .I(Decode1448_inst0_I),
    .O(Decode1448_inst0_O)
);
assign Decode1458_inst0_I = I;
Decode1458 Decode1458_inst0 (
    .I(Decode1458_inst0_I),
    .O(Decode1458_inst0_O)
);
assign Decode1468_inst0_I = I;
Decode1468 Decode1468_inst0 (
    .I(Decode1468_inst0_I),
    .O(Decode1468_inst0_O)
);
assign Decode1478_inst0_I = I;
Decode1478 Decode1478_inst0 (
    .I(Decode1478_inst0_I),
    .O(Decode1478_inst0_O)
);
assign Decode1488_inst0_I = I;
Decode1488 Decode1488_inst0 (
    .I(Decode1488_inst0_I),
    .O(Decode1488_inst0_O)
);
assign Decode148_inst0_I = I;
Decode148 Decode148_inst0 (
    .I(Decode148_inst0_I),
    .O(Decode148_inst0_O)
);
assign Decode1498_inst0_I = I;
Decode1498 Decode1498_inst0 (
    .I(Decode1498_inst0_I),
    .O(Decode1498_inst0_O)
);
assign Decode1508_inst0_I = I;
Decode1508 Decode1508_inst0 (
    .I(Decode1508_inst0_I),
    .O(Decode1508_inst0_O)
);
assign Decode1518_inst0_I = I;
Decode1518 Decode1518_inst0 (
    .I(Decode1518_inst0_I),
    .O(Decode1518_inst0_O)
);
assign Decode1528_inst0_I = I;
Decode1528 Decode1528_inst0 (
    .I(Decode1528_inst0_I),
    .O(Decode1528_inst0_O)
);
assign Decode1538_inst0_I = I;
Decode1538 Decode1538_inst0 (
    .I(Decode1538_inst0_I),
    .O(Decode1538_inst0_O)
);
assign Decode1548_inst0_I = I;
Decode1548 Decode1548_inst0 (
    .I(Decode1548_inst0_I),
    .O(Decode1548_inst0_O)
);
assign Decode1558_inst0_I = I;
Decode1558 Decode1558_inst0 (
    .I(Decode1558_inst0_I),
    .O(Decode1558_inst0_O)
);
assign Decode1568_inst0_I = I;
Decode1568 Decode1568_inst0 (
    .I(Decode1568_inst0_I),
    .O(Decode1568_inst0_O)
);
assign Decode1578_inst0_I = I;
Decode1578 Decode1578_inst0 (
    .I(Decode1578_inst0_I),
    .O(Decode1578_inst0_O)
);
assign Decode1588_inst0_I = I;
Decode1588 Decode1588_inst0 (
    .I(Decode1588_inst0_I),
    .O(Decode1588_inst0_O)
);
assign Decode158_inst0_I = I;
Decode158 Decode158_inst0 (
    .I(Decode158_inst0_I),
    .O(Decode158_inst0_O)
);
assign Decode1598_inst0_I = I;
Decode1598 Decode1598_inst0 (
    .I(Decode1598_inst0_I),
    .O(Decode1598_inst0_O)
);
assign Decode1608_inst0_I = I;
Decode1608 Decode1608_inst0 (
    .I(Decode1608_inst0_I),
    .O(Decode1608_inst0_O)
);
assign Decode1618_inst0_I = I;
Decode1618 Decode1618_inst0 (
    .I(Decode1618_inst0_I),
    .O(Decode1618_inst0_O)
);
assign Decode1628_inst0_I = I;
Decode1628 Decode1628_inst0 (
    .I(Decode1628_inst0_I),
    .O(Decode1628_inst0_O)
);
assign Decode1638_inst0_I = I;
Decode1638 Decode1638_inst0 (
    .I(Decode1638_inst0_I),
    .O(Decode1638_inst0_O)
);
assign Decode1648_inst0_I = I;
Decode1648 Decode1648_inst0 (
    .I(Decode1648_inst0_I),
    .O(Decode1648_inst0_O)
);
assign Decode1658_inst0_I = I;
Decode1658 Decode1658_inst0 (
    .I(Decode1658_inst0_I),
    .O(Decode1658_inst0_O)
);
assign Decode1668_inst0_I = I;
Decode1668 Decode1668_inst0 (
    .I(Decode1668_inst0_I),
    .O(Decode1668_inst0_O)
);
assign Decode1678_inst0_I = I;
Decode1678 Decode1678_inst0 (
    .I(Decode1678_inst0_I),
    .O(Decode1678_inst0_O)
);
assign Decode1688_inst0_I = I;
Decode1688 Decode1688_inst0 (
    .I(Decode1688_inst0_I),
    .O(Decode1688_inst0_O)
);
assign Decode168_inst0_I = I;
Decode168 Decode168_inst0 (
    .I(Decode168_inst0_I),
    .O(Decode168_inst0_O)
);
assign Decode1698_inst0_I = I;
Decode1698 Decode1698_inst0 (
    .I(Decode1698_inst0_I),
    .O(Decode1698_inst0_O)
);
assign Decode1708_inst0_I = I;
Decode1708 Decode1708_inst0 (
    .I(Decode1708_inst0_I),
    .O(Decode1708_inst0_O)
);
assign Decode1718_inst0_I = I;
Decode1718 Decode1718_inst0 (
    .I(Decode1718_inst0_I),
    .O(Decode1718_inst0_O)
);
assign Decode1728_inst0_I = I;
Decode1728 Decode1728_inst0 (
    .I(Decode1728_inst0_I),
    .O(Decode1728_inst0_O)
);
assign Decode1738_inst0_I = I;
Decode1738 Decode1738_inst0 (
    .I(Decode1738_inst0_I),
    .O(Decode1738_inst0_O)
);
assign Decode1748_inst0_I = I;
Decode1748 Decode1748_inst0 (
    .I(Decode1748_inst0_I),
    .O(Decode1748_inst0_O)
);
assign Decode1758_inst0_I = I;
Decode1758 Decode1758_inst0 (
    .I(Decode1758_inst0_I),
    .O(Decode1758_inst0_O)
);
assign Decode1768_inst0_I = I;
Decode1768 Decode1768_inst0 (
    .I(Decode1768_inst0_I),
    .O(Decode1768_inst0_O)
);
assign Decode1778_inst0_I = I;
Decode1778 Decode1778_inst0 (
    .I(Decode1778_inst0_I),
    .O(Decode1778_inst0_O)
);
assign Decode1788_inst0_I = I;
Decode1788 Decode1788_inst0 (
    .I(Decode1788_inst0_I),
    .O(Decode1788_inst0_O)
);
assign Decode178_inst0_I = I;
Decode178 Decode178_inst0 (
    .I(Decode178_inst0_I),
    .O(Decode178_inst0_O)
);
assign Decode1798_inst0_I = I;
Decode1798 Decode1798_inst0 (
    .I(Decode1798_inst0_I),
    .O(Decode1798_inst0_O)
);
assign Decode1808_inst0_I = I;
Decode1808 Decode1808_inst0 (
    .I(Decode1808_inst0_I),
    .O(Decode1808_inst0_O)
);
assign Decode1818_inst0_I = I;
Decode1818 Decode1818_inst0 (
    .I(Decode1818_inst0_I),
    .O(Decode1818_inst0_O)
);
assign Decode1828_inst0_I = I;
Decode1828 Decode1828_inst0 (
    .I(Decode1828_inst0_I),
    .O(Decode1828_inst0_O)
);
assign Decode1838_inst0_I = I;
Decode1838 Decode1838_inst0 (
    .I(Decode1838_inst0_I),
    .O(Decode1838_inst0_O)
);
assign Decode1848_inst0_I = I;
Decode1848 Decode1848_inst0 (
    .I(Decode1848_inst0_I),
    .O(Decode1848_inst0_O)
);
assign Decode1858_inst0_I = I;
Decode1858 Decode1858_inst0 (
    .I(Decode1858_inst0_I),
    .O(Decode1858_inst0_O)
);
assign Decode1868_inst0_I = I;
Decode1868 Decode1868_inst0 (
    .I(Decode1868_inst0_I),
    .O(Decode1868_inst0_O)
);
assign Decode1878_inst0_I = I;
Decode1878 Decode1878_inst0 (
    .I(Decode1878_inst0_I),
    .O(Decode1878_inst0_O)
);
assign Decode1888_inst0_I = I;
Decode1888 Decode1888_inst0 (
    .I(Decode1888_inst0_I),
    .O(Decode1888_inst0_O)
);
assign Decode188_inst0_I = I;
Decode188 Decode188_inst0 (
    .I(Decode188_inst0_I),
    .O(Decode188_inst0_O)
);
assign Decode1898_inst0_I = I;
Decode1898 Decode1898_inst0 (
    .I(Decode1898_inst0_I),
    .O(Decode1898_inst0_O)
);
assign Decode18_inst0_I = I;
Decode18 Decode18_inst0 (
    .I(Decode18_inst0_I),
    .O(Decode18_inst0_O)
);
assign Decode1908_inst0_I = I;
Decode1908 Decode1908_inst0 (
    .I(Decode1908_inst0_I),
    .O(Decode1908_inst0_O)
);
assign Decode1918_inst0_I = I;
Decode1918 Decode1918_inst0 (
    .I(Decode1918_inst0_I),
    .O(Decode1918_inst0_O)
);
assign Decode1928_inst0_I = I;
Decode1928 Decode1928_inst0 (
    .I(Decode1928_inst0_I),
    .O(Decode1928_inst0_O)
);
assign Decode1938_inst0_I = I;
Decode1938 Decode1938_inst0 (
    .I(Decode1938_inst0_I),
    .O(Decode1938_inst0_O)
);
assign Decode1948_inst0_I = I;
Decode1948 Decode1948_inst0 (
    .I(Decode1948_inst0_I),
    .O(Decode1948_inst0_O)
);
assign Decode1958_inst0_I = I;
Decode1958 Decode1958_inst0 (
    .I(Decode1958_inst0_I),
    .O(Decode1958_inst0_O)
);
assign Decode1968_inst0_I = I;
Decode1968 Decode1968_inst0 (
    .I(Decode1968_inst0_I),
    .O(Decode1968_inst0_O)
);
assign Decode1978_inst0_I = I;
Decode1978 Decode1978_inst0 (
    .I(Decode1978_inst0_I),
    .O(Decode1978_inst0_O)
);
assign Decode1988_inst0_I = I;
Decode1988 Decode1988_inst0 (
    .I(Decode1988_inst0_I),
    .O(Decode1988_inst0_O)
);
assign Decode198_inst0_I = I;
Decode198 Decode198_inst0 (
    .I(Decode198_inst0_I),
    .O(Decode198_inst0_O)
);
assign Decode1998_inst0_I = I;
Decode1998 Decode1998_inst0 (
    .I(Decode1998_inst0_I),
    .O(Decode1998_inst0_O)
);
assign Decode2008_inst0_I = I;
Decode2008 Decode2008_inst0 (
    .I(Decode2008_inst0_I),
    .O(Decode2008_inst0_O)
);
assign Decode2018_inst0_I = I;
Decode2018 Decode2018_inst0 (
    .I(Decode2018_inst0_I),
    .O(Decode2018_inst0_O)
);
assign Decode2028_inst0_I = I;
Decode2028 Decode2028_inst0 (
    .I(Decode2028_inst0_I),
    .O(Decode2028_inst0_O)
);
assign Decode2038_inst0_I = I;
Decode2038 Decode2038_inst0 (
    .I(Decode2038_inst0_I),
    .O(Decode2038_inst0_O)
);
assign Decode2048_inst0_I = I;
Decode2048 Decode2048_inst0 (
    .I(Decode2048_inst0_I),
    .O(Decode2048_inst0_O)
);
assign Decode2058_inst0_I = I;
Decode2058 Decode2058_inst0 (
    .I(Decode2058_inst0_I),
    .O(Decode2058_inst0_O)
);
assign Decode2068_inst0_I = I;
Decode2068 Decode2068_inst0 (
    .I(Decode2068_inst0_I),
    .O(Decode2068_inst0_O)
);
assign Decode2078_inst0_I = I;
Decode2078 Decode2078_inst0 (
    .I(Decode2078_inst0_I),
    .O(Decode2078_inst0_O)
);
assign Decode2088_inst0_I = I;
Decode2088 Decode2088_inst0 (
    .I(Decode2088_inst0_I),
    .O(Decode2088_inst0_O)
);
assign Decode208_inst0_I = I;
Decode208 Decode208_inst0 (
    .I(Decode208_inst0_I),
    .O(Decode208_inst0_O)
);
assign Decode2098_inst0_I = I;
Decode2098 Decode2098_inst0 (
    .I(Decode2098_inst0_I),
    .O(Decode2098_inst0_O)
);
assign Decode2108_inst0_I = I;
Decode2108 Decode2108_inst0 (
    .I(Decode2108_inst0_I),
    .O(Decode2108_inst0_O)
);
assign Decode2118_inst0_I = I;
Decode2118 Decode2118_inst0 (
    .I(Decode2118_inst0_I),
    .O(Decode2118_inst0_O)
);
assign Decode2128_inst0_I = I;
Decode2128 Decode2128_inst0 (
    .I(Decode2128_inst0_I),
    .O(Decode2128_inst0_O)
);
assign Decode2138_inst0_I = I;
Decode2138 Decode2138_inst0 (
    .I(Decode2138_inst0_I),
    .O(Decode2138_inst0_O)
);
assign Decode2148_inst0_I = I;
Decode2148 Decode2148_inst0 (
    .I(Decode2148_inst0_I),
    .O(Decode2148_inst0_O)
);
assign Decode2158_inst0_I = I;
Decode2158 Decode2158_inst0 (
    .I(Decode2158_inst0_I),
    .O(Decode2158_inst0_O)
);
assign Decode2168_inst0_I = I;
Decode2168 Decode2168_inst0 (
    .I(Decode2168_inst0_I),
    .O(Decode2168_inst0_O)
);
assign Decode2178_inst0_I = I;
Decode2178 Decode2178_inst0 (
    .I(Decode2178_inst0_I),
    .O(Decode2178_inst0_O)
);
assign Decode2188_inst0_I = I;
Decode2188 Decode2188_inst0 (
    .I(Decode2188_inst0_I),
    .O(Decode2188_inst0_O)
);
assign Decode218_inst0_I = I;
Decode218 Decode218_inst0 (
    .I(Decode218_inst0_I),
    .O(Decode218_inst0_O)
);
assign Decode2198_inst0_I = I;
Decode2198 Decode2198_inst0 (
    .I(Decode2198_inst0_I),
    .O(Decode2198_inst0_O)
);
assign Decode2208_inst0_I = I;
Decode2208 Decode2208_inst0 (
    .I(Decode2208_inst0_I),
    .O(Decode2208_inst0_O)
);
assign Decode2218_inst0_I = I;
Decode2218 Decode2218_inst0 (
    .I(Decode2218_inst0_I),
    .O(Decode2218_inst0_O)
);
assign Decode2228_inst0_I = I;
Decode2228 Decode2228_inst0 (
    .I(Decode2228_inst0_I),
    .O(Decode2228_inst0_O)
);
assign Decode2238_inst0_I = I;
Decode2238 Decode2238_inst0 (
    .I(Decode2238_inst0_I),
    .O(Decode2238_inst0_O)
);
assign Decode2248_inst0_I = I;
Decode2248 Decode2248_inst0 (
    .I(Decode2248_inst0_I),
    .O(Decode2248_inst0_O)
);
assign Decode2258_inst0_I = I;
Decode2258 Decode2258_inst0 (
    .I(Decode2258_inst0_I),
    .O(Decode2258_inst0_O)
);
assign Decode2268_inst0_I = I;
Decode2268 Decode2268_inst0 (
    .I(Decode2268_inst0_I),
    .O(Decode2268_inst0_O)
);
assign Decode2278_inst0_I = I;
Decode2278 Decode2278_inst0 (
    .I(Decode2278_inst0_I),
    .O(Decode2278_inst0_O)
);
assign Decode2288_inst0_I = I;
Decode2288 Decode2288_inst0 (
    .I(Decode2288_inst0_I),
    .O(Decode2288_inst0_O)
);
assign Decode228_inst0_I = I;
Decode228 Decode228_inst0 (
    .I(Decode228_inst0_I),
    .O(Decode228_inst0_O)
);
assign Decode2298_inst0_I = I;
Decode2298 Decode2298_inst0 (
    .I(Decode2298_inst0_I),
    .O(Decode2298_inst0_O)
);
assign Decode2308_inst0_I = I;
Decode2308 Decode2308_inst0 (
    .I(Decode2308_inst0_I),
    .O(Decode2308_inst0_O)
);
assign Decode2318_inst0_I = I;
Decode2318 Decode2318_inst0 (
    .I(Decode2318_inst0_I),
    .O(Decode2318_inst0_O)
);
assign Decode2328_inst0_I = I;
Decode2328 Decode2328_inst0 (
    .I(Decode2328_inst0_I),
    .O(Decode2328_inst0_O)
);
assign Decode2338_inst0_I = I;
Decode2338 Decode2338_inst0 (
    .I(Decode2338_inst0_I),
    .O(Decode2338_inst0_O)
);
assign Decode2348_inst0_I = I;
Decode2348 Decode2348_inst0 (
    .I(Decode2348_inst0_I),
    .O(Decode2348_inst0_O)
);
assign Decode2358_inst0_I = I;
Decode2358 Decode2358_inst0 (
    .I(Decode2358_inst0_I),
    .O(Decode2358_inst0_O)
);
assign Decode2368_inst0_I = I;
Decode2368 Decode2368_inst0 (
    .I(Decode2368_inst0_I),
    .O(Decode2368_inst0_O)
);
assign Decode2378_inst0_I = I;
Decode2378 Decode2378_inst0 (
    .I(Decode2378_inst0_I),
    .O(Decode2378_inst0_O)
);
assign Decode2388_inst0_I = I;
Decode2388 Decode2388_inst0 (
    .I(Decode2388_inst0_I),
    .O(Decode2388_inst0_O)
);
assign Decode238_inst0_I = I;
Decode238 Decode238_inst0 (
    .I(Decode238_inst0_I),
    .O(Decode238_inst0_O)
);
assign Decode2398_inst0_I = I;
Decode2398 Decode2398_inst0 (
    .I(Decode2398_inst0_I),
    .O(Decode2398_inst0_O)
);
assign Decode2408_inst0_I = I;
Decode2408 Decode2408_inst0 (
    .I(Decode2408_inst0_I),
    .O(Decode2408_inst0_O)
);
assign Decode2418_inst0_I = I;
Decode2418 Decode2418_inst0 (
    .I(Decode2418_inst0_I),
    .O(Decode2418_inst0_O)
);
assign Decode2428_inst0_I = I;
Decode2428 Decode2428_inst0 (
    .I(Decode2428_inst0_I),
    .O(Decode2428_inst0_O)
);
assign Decode2438_inst0_I = I;
Decode2438 Decode2438_inst0 (
    .I(Decode2438_inst0_I),
    .O(Decode2438_inst0_O)
);
assign Decode2448_inst0_I = I;
Decode2448 Decode2448_inst0 (
    .I(Decode2448_inst0_I),
    .O(Decode2448_inst0_O)
);
assign Decode2458_inst0_I = I;
Decode2458 Decode2458_inst0 (
    .I(Decode2458_inst0_I),
    .O(Decode2458_inst0_O)
);
assign Decode2468_inst0_I = I;
Decode2468 Decode2468_inst0 (
    .I(Decode2468_inst0_I),
    .O(Decode2468_inst0_O)
);
assign Decode2478_inst0_I = I;
Decode2478 Decode2478_inst0 (
    .I(Decode2478_inst0_I),
    .O(Decode2478_inst0_O)
);
assign Decode2488_inst0_I = I;
Decode2488 Decode2488_inst0 (
    .I(Decode2488_inst0_I),
    .O(Decode2488_inst0_O)
);
assign Decode248_inst0_I = I;
Decode248 Decode248_inst0 (
    .I(Decode248_inst0_I),
    .O(Decode248_inst0_O)
);
assign Decode2498_inst0_I = I;
Decode2498 Decode2498_inst0 (
    .I(Decode2498_inst0_I),
    .O(Decode2498_inst0_O)
);
assign Decode2508_inst0_I = I;
Decode2508 Decode2508_inst0 (
    .I(Decode2508_inst0_I),
    .O(Decode2508_inst0_O)
);
assign Decode2518_inst0_I = I;
Decode2518 Decode2518_inst0 (
    .I(Decode2518_inst0_I),
    .O(Decode2518_inst0_O)
);
assign Decode2528_inst0_I = I;
Decode2528 Decode2528_inst0 (
    .I(Decode2528_inst0_I),
    .O(Decode2528_inst0_O)
);
assign Decode2538_inst0_I = I;
Decode2538 Decode2538_inst0 (
    .I(Decode2538_inst0_I),
    .O(Decode2538_inst0_O)
);
assign Decode2548_inst0_I = I;
Decode2548 Decode2548_inst0 (
    .I(Decode2548_inst0_I),
    .O(Decode2548_inst0_O)
);
assign Decode2558_inst0_I = I;
Decode2558 Decode2558_inst0 (
    .I(Decode2558_inst0_I),
    .O(Decode2558_inst0_O)
);
assign Decode258_inst0_I = I;
Decode258 Decode258_inst0 (
    .I(Decode258_inst0_I),
    .O(Decode258_inst0_O)
);
assign Decode268_inst0_I = I;
Decode268 Decode268_inst0 (
    .I(Decode268_inst0_I),
    .O(Decode268_inst0_O)
);
assign Decode278_inst0_I = I;
Decode278 Decode278_inst0 (
    .I(Decode278_inst0_I),
    .O(Decode278_inst0_O)
);
assign Decode288_inst0_I = I;
Decode288 Decode288_inst0 (
    .I(Decode288_inst0_I),
    .O(Decode288_inst0_O)
);
assign Decode28_inst0_I = I;
Decode28 Decode28_inst0 (
    .I(Decode28_inst0_I),
    .O(Decode28_inst0_O)
);
assign Decode298_inst0_I = I;
Decode298 Decode298_inst0 (
    .I(Decode298_inst0_I),
    .O(Decode298_inst0_O)
);
assign Decode308_inst0_I = I;
Decode308 Decode308_inst0 (
    .I(Decode308_inst0_I),
    .O(Decode308_inst0_O)
);
assign Decode318_inst0_I = I;
Decode318 Decode318_inst0 (
    .I(Decode318_inst0_I),
    .O(Decode318_inst0_O)
);
assign Decode328_inst0_I = I;
Decode328 Decode328_inst0 (
    .I(Decode328_inst0_I),
    .O(Decode328_inst0_O)
);
assign Decode338_inst0_I = I;
Decode338 Decode338_inst0 (
    .I(Decode338_inst0_I),
    .O(Decode338_inst0_O)
);
assign Decode348_inst0_I = I;
Decode348 Decode348_inst0 (
    .I(Decode348_inst0_I),
    .O(Decode348_inst0_O)
);
assign Decode358_inst0_I = I;
Decode358 Decode358_inst0 (
    .I(Decode358_inst0_I),
    .O(Decode358_inst0_O)
);
assign Decode368_inst0_I = I;
Decode368 Decode368_inst0 (
    .I(Decode368_inst0_I),
    .O(Decode368_inst0_O)
);
assign Decode378_inst0_I = I;
Decode378 Decode378_inst0 (
    .I(Decode378_inst0_I),
    .O(Decode378_inst0_O)
);
assign Decode388_inst0_I = I;
Decode388 Decode388_inst0 (
    .I(Decode388_inst0_I),
    .O(Decode388_inst0_O)
);
assign Decode38_inst0_I = I;
Decode38 Decode38_inst0 (
    .I(Decode38_inst0_I),
    .O(Decode38_inst0_O)
);
assign Decode398_inst0_I = I;
Decode398 Decode398_inst0 (
    .I(Decode398_inst0_I),
    .O(Decode398_inst0_O)
);
assign Decode408_inst0_I = I;
Decode408 Decode408_inst0 (
    .I(Decode408_inst0_I),
    .O(Decode408_inst0_O)
);
assign Decode418_inst0_I = I;
Decode418 Decode418_inst0 (
    .I(Decode418_inst0_I),
    .O(Decode418_inst0_O)
);
assign Decode428_inst0_I = I;
Decode428 Decode428_inst0 (
    .I(Decode428_inst0_I),
    .O(Decode428_inst0_O)
);
assign Decode438_inst0_I = I;
Decode438 Decode438_inst0 (
    .I(Decode438_inst0_I),
    .O(Decode438_inst0_O)
);
assign Decode448_inst0_I = I;
Decode448 Decode448_inst0 (
    .I(Decode448_inst0_I),
    .O(Decode448_inst0_O)
);
assign Decode458_inst0_I = I;
Decode458 Decode458_inst0 (
    .I(Decode458_inst0_I),
    .O(Decode458_inst0_O)
);
assign Decode468_inst0_I = I;
Decode468 Decode468_inst0 (
    .I(Decode468_inst0_I),
    .O(Decode468_inst0_O)
);
assign Decode478_inst0_I = I;
Decode478 Decode478_inst0 (
    .I(Decode478_inst0_I),
    .O(Decode478_inst0_O)
);
assign Decode488_inst0_I = I;
Decode488 Decode488_inst0 (
    .I(Decode488_inst0_I),
    .O(Decode488_inst0_O)
);
assign Decode48_inst0_I = I;
Decode48 Decode48_inst0 (
    .I(Decode48_inst0_I),
    .O(Decode48_inst0_O)
);
assign Decode498_inst0_I = I;
Decode498 Decode498_inst0 (
    .I(Decode498_inst0_I),
    .O(Decode498_inst0_O)
);
assign Decode508_inst0_I = I;
Decode508 Decode508_inst0 (
    .I(Decode508_inst0_I),
    .O(Decode508_inst0_O)
);
assign Decode518_inst0_I = I;
Decode518 Decode518_inst0 (
    .I(Decode518_inst0_I),
    .O(Decode518_inst0_O)
);
assign Decode528_inst0_I = I;
Decode528 Decode528_inst0 (
    .I(Decode528_inst0_I),
    .O(Decode528_inst0_O)
);
assign Decode538_inst0_I = I;
Decode538 Decode538_inst0 (
    .I(Decode538_inst0_I),
    .O(Decode538_inst0_O)
);
assign Decode548_inst0_I = I;
Decode548 Decode548_inst0 (
    .I(Decode548_inst0_I),
    .O(Decode548_inst0_O)
);
assign Decode558_inst0_I = I;
Decode558 Decode558_inst0 (
    .I(Decode558_inst0_I),
    .O(Decode558_inst0_O)
);
assign Decode568_inst0_I = I;
Decode568 Decode568_inst0 (
    .I(Decode568_inst0_I),
    .O(Decode568_inst0_O)
);
assign Decode578_inst0_I = I;
Decode578 Decode578_inst0 (
    .I(Decode578_inst0_I),
    .O(Decode578_inst0_O)
);
assign Decode588_inst0_I = I;
Decode588 Decode588_inst0 (
    .I(Decode588_inst0_I),
    .O(Decode588_inst0_O)
);
assign Decode58_inst0_I = I;
Decode58 Decode58_inst0 (
    .I(Decode58_inst0_I),
    .O(Decode58_inst0_O)
);
assign Decode598_inst0_I = I;
Decode598 Decode598_inst0 (
    .I(Decode598_inst0_I),
    .O(Decode598_inst0_O)
);
assign Decode608_inst0_I = I;
Decode608 Decode608_inst0 (
    .I(Decode608_inst0_I),
    .O(Decode608_inst0_O)
);
assign Decode618_inst0_I = I;
Decode618 Decode618_inst0 (
    .I(Decode618_inst0_I),
    .O(Decode618_inst0_O)
);
assign Decode628_inst0_I = I;
Decode628 Decode628_inst0 (
    .I(Decode628_inst0_I),
    .O(Decode628_inst0_O)
);
assign Decode638_inst0_I = I;
Decode638 Decode638_inst0 (
    .I(Decode638_inst0_I),
    .O(Decode638_inst0_O)
);
assign Decode648_inst0_I = I;
Decode648 Decode648_inst0 (
    .I(Decode648_inst0_I),
    .O(Decode648_inst0_O)
);
assign Decode658_inst0_I = I;
Decode658 Decode658_inst0 (
    .I(Decode658_inst0_I),
    .O(Decode658_inst0_O)
);
assign Decode668_inst0_I = I;
Decode668 Decode668_inst0 (
    .I(Decode668_inst0_I),
    .O(Decode668_inst0_O)
);
assign Decode678_inst0_I = I;
Decode678 Decode678_inst0 (
    .I(Decode678_inst0_I),
    .O(Decode678_inst0_O)
);
assign Decode688_inst0_I = I;
Decode688 Decode688_inst0 (
    .I(Decode688_inst0_I),
    .O(Decode688_inst0_O)
);
assign Decode68_inst0_I = I;
Decode68 Decode68_inst0 (
    .I(Decode68_inst0_I),
    .O(Decode68_inst0_O)
);
assign Decode698_inst0_I = I;
Decode698 Decode698_inst0 (
    .I(Decode698_inst0_I),
    .O(Decode698_inst0_O)
);
assign Decode708_inst0_I = I;
Decode708 Decode708_inst0 (
    .I(Decode708_inst0_I),
    .O(Decode708_inst0_O)
);
assign Decode718_inst0_I = I;
Decode718 Decode718_inst0 (
    .I(Decode718_inst0_I),
    .O(Decode718_inst0_O)
);
assign Decode728_inst0_I = I;
Decode728 Decode728_inst0 (
    .I(Decode728_inst0_I),
    .O(Decode728_inst0_O)
);
assign Decode738_inst0_I = I;
Decode738 Decode738_inst0 (
    .I(Decode738_inst0_I),
    .O(Decode738_inst0_O)
);
assign Decode748_inst0_I = I;
Decode748 Decode748_inst0 (
    .I(Decode748_inst0_I),
    .O(Decode748_inst0_O)
);
assign Decode758_inst0_I = I;
Decode758 Decode758_inst0 (
    .I(Decode758_inst0_I),
    .O(Decode758_inst0_O)
);
assign Decode768_inst0_I = I;
Decode768 Decode768_inst0 (
    .I(Decode768_inst0_I),
    .O(Decode768_inst0_O)
);
assign Decode778_inst0_I = I;
Decode778 Decode778_inst0 (
    .I(Decode778_inst0_I),
    .O(Decode778_inst0_O)
);
assign Decode788_inst0_I = I;
Decode788 Decode788_inst0 (
    .I(Decode788_inst0_I),
    .O(Decode788_inst0_O)
);
assign Decode78_inst0_I = I;
Decode78 Decode78_inst0 (
    .I(Decode78_inst0_I),
    .O(Decode78_inst0_O)
);
assign Decode798_inst0_I = I;
Decode798 Decode798_inst0 (
    .I(Decode798_inst0_I),
    .O(Decode798_inst0_O)
);
assign Decode808_inst0_I = I;
Decode808 Decode808_inst0 (
    .I(Decode808_inst0_I),
    .O(Decode808_inst0_O)
);
assign Decode818_inst0_I = I;
Decode818 Decode818_inst0 (
    .I(Decode818_inst0_I),
    .O(Decode818_inst0_O)
);
assign Decode828_inst0_I = I;
Decode828 Decode828_inst0 (
    .I(Decode828_inst0_I),
    .O(Decode828_inst0_O)
);
assign Decode838_inst0_I = I;
Decode838 Decode838_inst0 (
    .I(Decode838_inst0_I),
    .O(Decode838_inst0_O)
);
assign Decode848_inst0_I = I;
Decode848 Decode848_inst0 (
    .I(Decode848_inst0_I),
    .O(Decode848_inst0_O)
);
assign Decode858_inst0_I = I;
Decode858 Decode858_inst0 (
    .I(Decode858_inst0_I),
    .O(Decode858_inst0_O)
);
assign Decode868_inst0_I = I;
Decode868 Decode868_inst0 (
    .I(Decode868_inst0_I),
    .O(Decode868_inst0_O)
);
assign Decode878_inst0_I = I;
Decode878 Decode878_inst0 (
    .I(Decode878_inst0_I),
    .O(Decode878_inst0_O)
);
assign Decode888_inst0_I = I;
Decode888 Decode888_inst0 (
    .I(Decode888_inst0_I),
    .O(Decode888_inst0_O)
);
assign Decode88_inst0_I = I;
Decode88 Decode88_inst0 (
    .I(Decode88_inst0_I),
    .O(Decode88_inst0_O)
);
assign Decode898_inst0_I = I;
Decode898 Decode898_inst0 (
    .I(Decode898_inst0_I),
    .O(Decode898_inst0_O)
);
assign Decode908_inst0_I = I;
Decode908 Decode908_inst0 (
    .I(Decode908_inst0_I),
    .O(Decode908_inst0_O)
);
assign Decode918_inst0_I = I;
Decode918 Decode918_inst0 (
    .I(Decode918_inst0_I),
    .O(Decode918_inst0_O)
);
assign Decode928_inst0_I = I;
Decode928 Decode928_inst0 (
    .I(Decode928_inst0_I),
    .O(Decode928_inst0_O)
);
assign Decode938_inst0_I = I;
Decode938 Decode938_inst0 (
    .I(Decode938_inst0_I),
    .O(Decode938_inst0_O)
);
assign Decode948_inst0_I = I;
Decode948 Decode948_inst0 (
    .I(Decode948_inst0_I),
    .O(Decode948_inst0_O)
);
assign Decode958_inst0_I = I;
Decode958 Decode958_inst0 (
    .I(Decode958_inst0_I),
    .O(Decode958_inst0_O)
);
assign Decode968_inst0_I = I;
Decode968 Decode968_inst0 (
    .I(Decode968_inst0_I),
    .O(Decode968_inst0_O)
);
assign Decode978_inst0_I = I;
Decode978 Decode978_inst0 (
    .I(Decode978_inst0_I),
    .O(Decode978_inst0_O)
);
assign Decode988_inst0_I = I;
Decode988 Decode988_inst0 (
    .I(Decode988_inst0_I),
    .O(Decode988_inst0_O)
);
assign Decode98_inst0_I = I;
Decode98 Decode98_inst0 (
    .I(Decode98_inst0_I),
    .O(Decode98_inst0_O)
);
assign Decode998_inst0_I = I;
Decode998 Decode998_inst0 (
    .I(Decode998_inst0_I),
    .O(Decode998_inst0_O)
);
assign O = {Decode2558_inst0_O,Decode2548_inst0_O,Decode2538_inst0_O,Decode2528_inst0_O,Decode2518_inst0_O,Decode2508_inst0_O,Decode2498_inst0_O,Decode2488_inst0_O,Decode2478_inst0_O,Decode2468_inst0_O,Decode2458_inst0_O,Decode2448_inst0_O,Decode2438_inst0_O,Decode2428_inst0_O,Decode2418_inst0_O,Decode2408_inst0_O,Decode2398_inst0_O,Decode2388_inst0_O,Decode2378_inst0_O,Decode2368_inst0_O,Decode2358_inst0_O,Decode2348_inst0_O,Decode2338_inst0_O,Decode2328_inst0_O,Decode2318_inst0_O,Decode2308_inst0_O,Decode2298_inst0_O,Decode2288_inst0_O,Decode2278_inst0_O,Decode2268_inst0_O,Decode2258_inst0_O,Decode2248_inst0_O,Decode2238_inst0_O,Decode2228_inst0_O,Decode2218_inst0_O,Decode2208_inst0_O,Decode2198_inst0_O,Decode2188_inst0_O,Decode2178_inst0_O,Decode2168_inst0_O,Decode2158_inst0_O,Decode2148_inst0_O,Decode2138_inst0_O,Decode2128_inst0_O,Decode2118_inst0_O,Decode2108_inst0_O,Decode2098_inst0_O,Decode2088_inst0_O,Decode2078_inst0_O,Decode2068_inst0_O,Decode2058_inst0_O,Decode2048_inst0_O,Decode2038_inst0_O,Decode2028_inst0_O,Decode2018_inst0_O,Decode2008_inst0_O,Decode1998_inst0_O,Decode1988_inst0_O,Decode1978_inst0_O,Decode1968_inst0_O,Decode1958_inst0_O,Decode1948_inst0_O,Decode1938_inst0_O,Decode1928_inst0_O,Decode1918_inst0_O,Decode1908_inst0_O,Decode1898_inst0_O,Decode1888_inst0_O,Decode1878_inst0_O,Decode1868_inst0_O,Decode1858_inst0_O,Decode1848_inst0_O,Decode1838_inst0_O,Decode1828_inst0_O,Decode1818_inst0_O,Decode1808_inst0_O,Decode1798_inst0_O,Decode1788_inst0_O,Decode1778_inst0_O,Decode1768_inst0_O,Decode1758_inst0_O,Decode1748_inst0_O,Decode1738_inst0_O,Decode1728_inst0_O,Decode1718_inst0_O,Decode1708_inst0_O,Decode1698_inst0_O,Decode1688_inst0_O,Decode1678_inst0_O,Decode1668_inst0_O,Decode1658_inst0_O,Decode1648_inst0_O,Decode1638_inst0_O,Decode1628_inst0_O,Decode1618_inst0_O,Decode1608_inst0_O,Decode1598_inst0_O,Decode1588_inst0_O,Decode1578_inst0_O,Decode1568_inst0_O,Decode1558_inst0_O,Decode1548_inst0_O,Decode1538_inst0_O,Decode1528_inst0_O,Decode1518_inst0_O,Decode1508_inst0_O,Decode1498_inst0_O,Decode1488_inst0_O,Decode1478_inst0_O,Decode1468_inst0_O,Decode1458_inst0_O,Decode1448_inst0_O,Decode1438_inst0_O,Decode1428_inst0_O,Decode1418_inst0_O,Decode1408_inst0_O,Decode1398_inst0_O,Decode1388_inst0_O,Decode1378_inst0_O,Decode1368_inst0_O,Decode1358_inst0_O,Decode1348_inst0_O,Decode1338_inst0_O,Decode1328_inst0_O,Decode1318_inst0_O,Decode1308_inst0_O,Decode1298_inst0_O,Decode1288_inst0_O,Decode1278_inst0_O,Decode1268_inst0_O,Decode1258_inst0_O,Decode1248_inst0_O,Decode1238_inst0_O,Decode1228_inst0_O,Decode1218_inst0_O,Decode1208_inst0_O,Decode1198_inst0_O,Decode1188_inst0_O,Decode1178_inst0_O,Decode1168_inst0_O,Decode1158_inst0_O,Decode1148_inst0_O,Decode1138_inst0_O,Decode1128_inst0_O,Decode1118_inst0_O,Decode1108_inst0_O,Decode1098_inst0_O,Decode1088_inst0_O,Decode1078_inst0_O,Decode1068_inst0_O,Decode1058_inst0_O,Decode1048_inst0_O,Decode1038_inst0_O,Decode1028_inst0_O,Decode1018_inst0_O,Decode1008_inst0_O,Decode998_inst0_O,Decode988_inst0_O,Decode978_inst0_O,Decode968_inst0_O,Decode958_inst0_O,Decode948_inst0_O,Decode938_inst0_O,Decode928_inst0_O,Decode918_inst0_O,Decode908_inst0_O,Decode898_inst0_O,Decode888_inst0_O,Decode878_inst0_O,Decode868_inst0_O,Decode858_inst0_O,Decode848_inst0_O,Decode838_inst0_O,Decode828_inst0_O,Decode818_inst0_O,Decode808_inst0_O,Decode798_inst0_O,Decode788_inst0_O,Decode778_inst0_O,Decode768_inst0_O,Decode758_inst0_O,Decode748_inst0_O,Decode738_inst0_O,Decode728_inst0_O,Decode718_inst0_O,Decode708_inst0_O,Decode698_inst0_O,Decode688_inst0_O,Decode678_inst0_O,Decode668_inst0_O,Decode658_inst0_O,Decode648_inst0_O,Decode638_inst0_O,Decode628_inst0_O,Decode618_inst0_O,Decode608_inst0_O,Decode598_inst0_O,Decode588_inst0_O,Decode578_inst0_O,Decode568_inst0_O,Decode558_inst0_O,Decode548_inst0_O,Decode538_inst0_O,Decode528_inst0_O,Decode518_inst0_O,Decode508_inst0_O,Decode498_inst0_O,Decode488_inst0_O,Decode478_inst0_O,Decode468_inst0_O,Decode458_inst0_O,Decode448_inst0_O,Decode438_inst0_O,Decode428_inst0_O,Decode418_inst0_O,Decode408_inst0_O,Decode398_inst0_O,Decode388_inst0_O,Decode378_inst0_O,Decode368_inst0_O,Decode358_inst0_O,Decode348_inst0_O,Decode338_inst0_O,Decode328_inst0_O,Decode318_inst0_O,Decode308_inst0_O,Decode298_inst0_O,Decode288_inst0_O,Decode278_inst0_O,Decode268_inst0_O,Decode258_inst0_O,Decode248_inst0_O,Decode238_inst0_O,Decode228_inst0_O,Decode218_inst0_O,Decode208_inst0_O,Decode198_inst0_O,Decode188_inst0_O,Decode178_inst0_O,Decode168_inst0_O,Decode158_inst0_O,Decode148_inst0_O,Decode138_inst0_O,Decode128_inst0_O,Decode118_inst0_O,Decode108_inst0_O,Decode98_inst0_O,Decode88_inst0_O,Decode78_inst0_O,Decode68_inst0_O,Decode58_inst0_O,Decode48_inst0_O,Decode38_inst0_O,Decode28_inst0_O,Decode18_inst0_O,Decode08_inst0_O};
endmodule

