module Sub8_cin_cout (input [7:0] I0, input [7:0] I1, input  CIN, output [7:0] O, output  COUT);
wire  LUT6_2_inst0_O5;
wire  LUT6_2_inst0_O6;
wire  MUXCY_inst0_O;
wire  XORCY_inst0_O;
wire  LUT6_2_inst1_O5;
wire  LUT6_2_inst1_O6;
wire  MUXCY_inst1_O;
wire  XORCY_inst1_O;
wire  LUT6_2_inst2_O5;
wire  LUT6_2_inst2_O6;
wire  MUXCY_inst2_O;
wire  XORCY_inst2_O;
wire  LUT6_2_inst3_O5;
wire  LUT6_2_inst3_O6;
wire  MUXCY_inst3_O;
wire  XORCY_inst3_O;
wire  LUT6_2_inst4_O5;
wire  LUT6_2_inst4_O6;
wire  MUXCY_inst4_O;
wire  XORCY_inst4_O;
wire  LUT6_2_inst5_O5;
wire  LUT6_2_inst5_O6;
wire  MUXCY_inst5_O;
wire  XORCY_inst5_O;
wire  LUT6_2_inst6_O5;
wire  LUT6_2_inst6_O6;
wire  MUXCY_inst6_O;
wire  XORCY_inst6_O;
wire  LUT6_2_inst7_O5;
wire  LUT6_2_inst7_O6;
wire  MUXCY_inst7_O;
wire  XORCY_inst7_O;
wire  LUT1_inst0_O;
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst0 (.I0(I0[0]), .I1(I1[0]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst0_O5), .O6(LUT6_2_inst0_O6));
MUXCY MUXCY_inst0 (.DI(LUT6_2_inst0_O5), .CI(LUT1_inst0_O), .S(LUT6_2_inst0_O6), .O(MUXCY_inst0_O));
XORCY XORCY_inst0 (.LI(LUT6_2_inst0_O6), .CI(LUT1_inst0_O), .O(XORCY_inst0_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst1 (.I0(I0[1]), .I1(I1[1]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst1_O5), .O6(LUT6_2_inst1_O6));
MUXCY MUXCY_inst1 (.DI(LUT6_2_inst1_O5), .CI(MUXCY_inst0_O), .S(LUT6_2_inst1_O6), .O(MUXCY_inst1_O));
XORCY XORCY_inst1 (.LI(LUT6_2_inst1_O6), .CI(MUXCY_inst0_O), .O(XORCY_inst1_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst2 (.I0(I0[2]), .I1(I1[2]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst2_O5), .O6(LUT6_2_inst2_O6));
MUXCY MUXCY_inst2 (.DI(LUT6_2_inst2_O5), .CI(MUXCY_inst1_O), .S(LUT6_2_inst2_O6), .O(MUXCY_inst2_O));
XORCY XORCY_inst2 (.LI(LUT6_2_inst2_O6), .CI(MUXCY_inst1_O), .O(XORCY_inst2_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst3 (.I0(I0[3]), .I1(I1[3]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst3_O5), .O6(LUT6_2_inst3_O6));
MUXCY MUXCY_inst3 (.DI(LUT6_2_inst3_O5), .CI(MUXCY_inst2_O), .S(LUT6_2_inst3_O6), .O(MUXCY_inst3_O));
XORCY XORCY_inst3 (.LI(LUT6_2_inst3_O6), .CI(MUXCY_inst2_O), .O(XORCY_inst3_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst4 (.I0(I0[4]), .I1(I1[4]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst4_O5), .O6(LUT6_2_inst4_O6));
MUXCY MUXCY_inst4 (.DI(LUT6_2_inst4_O5), .CI(MUXCY_inst3_O), .S(LUT6_2_inst4_O6), .O(MUXCY_inst4_O));
XORCY XORCY_inst4 (.LI(LUT6_2_inst4_O6), .CI(MUXCY_inst3_O), .O(XORCY_inst4_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst5 (.I0(I0[5]), .I1(I1[5]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst5_O5), .O6(LUT6_2_inst5_O6));
MUXCY MUXCY_inst5 (.DI(LUT6_2_inst5_O5), .CI(MUXCY_inst4_O), .S(LUT6_2_inst5_O6), .O(MUXCY_inst5_O));
XORCY XORCY_inst5 (.LI(LUT6_2_inst5_O6), .CI(MUXCY_inst4_O), .O(XORCY_inst5_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst6 (.I0(I0[6]), .I1(I1[6]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst6_O5), .O6(LUT6_2_inst6_O6));
MUXCY MUXCY_inst6 (.DI(LUT6_2_inst6_O5), .CI(MUXCY_inst5_O), .S(LUT6_2_inst6_O6), .O(MUXCY_inst6_O));
XORCY XORCY_inst6 (.LI(LUT6_2_inst6_O6), .CI(MUXCY_inst5_O), .O(XORCY_inst6_O));
LUT6_2 #(.INIT(64'h99999999AAAAAAAA)) LUT6_2_inst7 (.I0(I0[7]), .I1(I1[7]), .I2(1'b0), .I3(1'b0), .I4(1'b0), .I5(1'b1), .O5(LUT6_2_inst7_O5), .O6(LUT6_2_inst7_O6));
MUXCY MUXCY_inst7 (.DI(LUT6_2_inst7_O5), .CI(MUXCY_inst6_O), .S(LUT6_2_inst7_O6), .O(MUXCY_inst7_O));
XORCY XORCY_inst7 (.LI(LUT6_2_inst7_O6), .CI(MUXCY_inst6_O), .O(XORCY_inst7_O));
LUT1 #(.INIT(2'h1)) LUT1_inst0 (.I0(CIN), .O(LUT1_inst0_O));
assign O = {XORCY_inst7_O,XORCY_inst6_O,XORCY_inst5_O,XORCY_inst4_O,XORCY_inst3_O,XORCY_inst2_O,XORCY_inst1_O,XORCY_inst0_O};
assign COUT = MUXCY_inst7_O;
endmodule

